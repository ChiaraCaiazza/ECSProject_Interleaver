------------------------------------------------------------------------------ -
--Interleaver - TestBench
--
--File name : interleaver_test-3.vhdl.vhdl
-- 
--Library : IEEE
--Author: Chiara Caiazza


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ieee.numeric_std.ALL;
 
ENTITY interleaver_test IS

END interleaver_test;

ARCHITECTURE interleaver_test_arch OF interleaver_test IS
	COMPONENT interleaver IS
		port(	clk : in std_logic;					--Processing clock
				reset : in  std_logic;				--Asynchronous active high reset
				bit_in : in std_logic;				--input bit
				bit_out : out std_logic				--outputbit
		);
	END COMPONENT interleaver;


	--CONSTANT
	CONSTANT clock_period : TIME := 200 ns;
	CONSTANT len : INTEGER := 2049;


	--INPUT SIGNALS
	SIGNAL clock : std_logic := '0';
	SIGNAL rst : std_logic := '1';
	SIGNAL bit_input : std_logic := '0';


	--OUTPUT SIGNALS
	SIGNAL bit_output : std_logic := 'Z';

	SIGNAL clock_cycle : INTEGER;
	SIGNAL testing: Boolean :=True;

	BEGIN
		I: interleaver PORT MAP(clk => clock, reset => rst, bit_in => bit_input, bit_out =>bit_output);

--Generates clk
		clock <=NOT clock AFTER clock_period/2 WHEN testing ELSE '0';

		--Runs simulation for len cycles
		proc_test: PROCESS(clock)
			VARIABLE count: INTEGER:= 0;
			BEGIN
				clock_cycle <= (count+1)/2;
				CASE count IS
					-- reset 
					WHEN	0	=>	rst<='1';

					-- starting input
					WHEN	1	=>	bit_input<='1';rst<='0';
					WHEN	2	=>	bit_input<='1';
					WHEN	3	=>	bit_input<='1';
					WHEN	4	=>	bit_input<='1';
					WHEN	5	=>	bit_input<='1';
					WHEN	6	=>	bit_input<='1';
					WHEN	7	=>	bit_input<='1';
					WHEN	8	=>	bit_input<='1';
					WHEN	9	=>	bit_input<='1';
					WHEN	10	=>	bit_input<='1';
					WHEN	11	=>	bit_input<='1';
					WHEN	12	=>	bit_input<='1';
					WHEN	13	=>	bit_input<='1';
					WHEN	14	=>	bit_input<='1';
					WHEN	15	=>	bit_input<='1';
					WHEN	16	=>	bit_input<='1';
					WHEN	17	=>	bit_input<='1';
					WHEN	18	=>	bit_input<='1';
					WHEN	19	=>	bit_input<='1';
					WHEN	20	=>	bit_input<='1';
					WHEN	21	=>	bit_input<='1';
					WHEN	22	=>	bit_input<='1';
					WHEN	23	=>	bit_input<='1';
					WHEN	24	=>	bit_input<='1';
					WHEN	25	=>	bit_input<='1';
					WHEN	26	=>	bit_input<='1';
					WHEN	27	=>	bit_input<='1';
					WHEN	28	=>	bit_input<='1';
					WHEN	29	=>	bit_input<='1';
					WHEN	30	=>	bit_input<='1';
					WHEN	31	=>	bit_input<='1';
					WHEN	32	=>	bit_input<='1';
					WHEN	33	=>	bit_input<='1';
					WHEN	34	=>	bit_input<='1';
					WHEN	35	=>	bit_input<='1';
					WHEN	36	=>	bit_input<='1';
					WHEN	37	=>	bit_input<='1';
					WHEN	38	=>	bit_input<='1';
					WHEN	39	=>	bit_input<='1';
					WHEN	40	=>	bit_input<='1';
					WHEN	41	=>	bit_input<='1';
					WHEN	42	=>	bit_input<='1';
					WHEN	43	=>	bit_input<='1';
					WHEN	44	=>	bit_input<='1';
					WHEN	45	=>	bit_input<='1';
					WHEN	46	=>	bit_input<='1';
					WHEN	47	=>	bit_input<='1';
					WHEN	48	=>	bit_input<='1';
					WHEN	49	=>	bit_input<='1';
					WHEN	50	=>	bit_input<='1';
					WHEN	51	=>	bit_input<='1';
					WHEN	52	=>	bit_input<='1';
					WHEN	53	=>	bit_input<='1';
					WHEN	54	=>	bit_input<='1';
					WHEN	55	=>	bit_input<='1';
					WHEN	56	=>	bit_input<='1';
					WHEN	57	=>	bit_input<='1';
					WHEN	58	=>	bit_input<='1';
					WHEN	59	=>	bit_input<='1';
					WHEN	60	=>	bit_input<='1';
					WHEN	61	=>	bit_input<='1';
					WHEN	62	=>	bit_input<='1';
					WHEN	63	=>	bit_input<='1';
					WHEN	64	=>	bit_input<='1';
					WHEN	65	=>	bit_input<='1';
					WHEN	66	=>	bit_input<='1';
					WHEN	67	=>	bit_input<='1';
					WHEN	68	=>	bit_input<='1';
					WHEN	69	=>	bit_input<='1';
					WHEN	70	=>	bit_input<='1';
					WHEN	71	=>	bit_input<='1';
					WHEN	72	=>	bit_input<='1';
					WHEN	73	=>	bit_input<='1';
					WHEN	74	=>	bit_input<='1';
					WHEN	75	=>	bit_input<='1';
					WHEN	76	=>	bit_input<='1';
					WHEN	77	=>	bit_input<='1';
					WHEN	78	=>	bit_input<='1';
					WHEN	79	=>	bit_input<='1';
					WHEN	80	=>	bit_input<='1';
					WHEN	81	=>	bit_input<='1';
					WHEN	82	=>	bit_input<='1';
					WHEN	83	=>	bit_input<='1';
					WHEN	84	=>	bit_input<='1';
					WHEN	85	=>	bit_input<='1';
					WHEN	86	=>	bit_input<='1';
					WHEN	87	=>	bit_input<='1';
					WHEN	88	=>	bit_input<='1';
					WHEN	89	=>	bit_input<='1';
					WHEN	90	=>	bit_input<='1';
					WHEN	91	=>	bit_input<='1';
					WHEN	92	=>	bit_input<='1';
					WHEN	93	=>	bit_input<='1';
					WHEN	94	=>	bit_input<='1';
					WHEN	95	=>	bit_input<='1';
					WHEN	96	=>	bit_input<='1';
					WHEN	97	=>	bit_input<='1';
					WHEN	98	=>	bit_input<='1';
					WHEN	99	=>	bit_input<='1';
					WHEN	100	=>	bit_input<='1';
					WHEN	101	=>	bit_input<='1';
					WHEN	102	=>	bit_input<='1';
					WHEN	103	=>	bit_input<='1';
					WHEN	104	=>	bit_input<='1';
					WHEN	105	=>	bit_input<='1';
					WHEN	106	=>	bit_input<='1';
					WHEN	107	=>	bit_input<='1';
					WHEN	108	=>	bit_input<='1';
					WHEN	109	=>	bit_input<='1';
					WHEN	110	=>	bit_input<='1';
					WHEN	111	=>	bit_input<='1';
					WHEN	112	=>	bit_input<='1';
					WHEN	113	=>	bit_input<='1';
					WHEN	114	=>	bit_input<='1';
					WHEN	115	=>	bit_input<='1';
					WHEN	116	=>	bit_input<='1';
					WHEN	117	=>	bit_input<='1';
					WHEN	118	=>	bit_input<='1';
					WHEN	119	=>	bit_input<='1';
					WHEN	120	=>	bit_input<='1';
					WHEN	121	=>	bit_input<='1';
					WHEN	122	=>	bit_input<='1';
					WHEN	123	=>	bit_input<='1';
					WHEN	124	=>	bit_input<='1';
					WHEN	125	=>	bit_input<='1';
					WHEN	126	=>	bit_input<='1';
					WHEN	127	=>	bit_input<='1';
					WHEN	128	=>	bit_input<='1';
					WHEN	129	=>	bit_input<='1';
					WHEN	130	=>	bit_input<='1';
					WHEN	131	=>	bit_input<='1';
					WHEN	132	=>	bit_input<='1';
					WHEN	133	=>	bit_input<='1';
					WHEN	134	=>	bit_input<='1';
					WHEN	135	=>	bit_input<='1';
					WHEN	136	=>	bit_input<='1';
					WHEN	137	=>	bit_input<='1';
					WHEN	138	=>	bit_input<='1';
					WHEN	139	=>	bit_input<='1';
					WHEN	140	=>	bit_input<='1';
					WHEN	141	=>	bit_input<='1';
					WHEN	142	=>	bit_input<='1';
					WHEN	143	=>	bit_input<='1';
					WHEN	144	=>	bit_input<='1';
					WHEN	145	=>	bit_input<='1';
					WHEN	146	=>	bit_input<='1';
					WHEN	147	=>	bit_input<='1';
					WHEN	148	=>	bit_input<='1';
					WHEN	149	=>	bit_input<='1';
					WHEN	150	=>	bit_input<='1';
					WHEN	151	=>	bit_input<='1';
					WHEN	152	=>	bit_input<='1';
					WHEN	153	=>	bit_input<='1';
					WHEN	154	=>	bit_input<='1';
					WHEN	155	=>	bit_input<='1';
					WHEN	156	=>	bit_input<='1';
					WHEN	157	=>	bit_input<='1';
					WHEN	158	=>	bit_input<='1';
					WHEN	159	=>	bit_input<='1';
					WHEN	160	=>	bit_input<='1';
					WHEN	161	=>	bit_input<='1';
					WHEN	162	=>	bit_input<='1';
					WHEN	163	=>	bit_input<='1';
					WHEN	164	=>	bit_input<='1';
					WHEN	165	=>	bit_input<='1';
					WHEN	166	=>	bit_input<='1';
					WHEN	167	=>	bit_input<='1';
					WHEN	168	=>	bit_input<='1';
					WHEN	169	=>	bit_input<='1';
					WHEN	170	=>	bit_input<='1';
					WHEN	171	=>	bit_input<='1';
					WHEN	172	=>	bit_input<='1';
					WHEN	173	=>	bit_input<='1';
					WHEN	174	=>	bit_input<='1';
					WHEN	175	=>	bit_input<='1';
					WHEN	176	=>	bit_input<='1';
					WHEN	177	=>	bit_input<='1';
					WHEN	178	=>	bit_input<='1';
					WHEN	179	=>	bit_input<='1';
					WHEN	180	=>	bit_input<='1';
					WHEN	181	=>	bit_input<='1';
					WHEN	182	=>	bit_input<='1';
					WHEN	183	=>	bit_input<='1';
					WHEN	184	=>	bit_input<='1';
					WHEN	185	=>	bit_input<='1';
					WHEN	186	=>	bit_input<='1';
					WHEN	187	=>	bit_input<='1';
					WHEN	188	=>	bit_input<='1';
					WHEN	189	=>	bit_input<='1';
					WHEN	190	=>	bit_input<='1';
					WHEN	191	=>	bit_input<='1';
					WHEN	192	=>	bit_input<='1';
					WHEN	193	=>	bit_input<='1';
					WHEN	194	=>	bit_input<='1';
					WHEN	195	=>	bit_input<='1';
					WHEN	196	=>	bit_input<='1';
					WHEN	197	=>	bit_input<='1';
					WHEN	198	=>	bit_input<='1';
					WHEN	199	=>	bit_input<='1';
					WHEN	200	=>	bit_input<='1';
					WHEN	201	=>	bit_input<='1';
					WHEN	202	=>	bit_input<='1';
					WHEN	203	=>	bit_input<='1';
					WHEN	204	=>	bit_input<='1';
					WHEN	205	=>	bit_input<='1';
					WHEN	206	=>	bit_input<='1';
					WHEN	207	=>	bit_input<='1';
					WHEN	208	=>	bit_input<='1';
					WHEN	209	=>	bit_input<='1';
					WHEN	210	=>	bit_input<='1';
					WHEN	211	=>	bit_input<='1';
					WHEN	212	=>	bit_input<='1';
					WHEN	213	=>	bit_input<='1';
					WHEN	214	=>	bit_input<='1';
					WHEN	215	=>	bit_input<='1';
					WHEN	216	=>	bit_input<='1';
					WHEN	217	=>	bit_input<='1';
					WHEN	218	=>	bit_input<='1';
					WHEN	219	=>	bit_input<='1';
					WHEN	220	=>	bit_input<='1';
					WHEN	221	=>	bit_input<='1';
					WHEN	222	=>	bit_input<='1';
					WHEN	223	=>	bit_input<='1';
					WHEN	224	=>	bit_input<='1';
					WHEN	225	=>	bit_input<='1';
					WHEN	226	=>	bit_input<='1';
					WHEN	227	=>	bit_input<='1';
					WHEN	228	=>	bit_input<='1';
					WHEN	229	=>	bit_input<='1';
					WHEN	230	=>	bit_input<='1';
					WHEN	231	=>	bit_input<='1';
					WHEN	232	=>	bit_input<='1';
					WHEN	233	=>	bit_input<='1';
					WHEN	234	=>	bit_input<='1';
					WHEN	235	=>	bit_input<='1';
					WHEN	236	=>	bit_input<='1';
					WHEN	237	=>	bit_input<='1';
					WHEN	238	=>	bit_input<='1';
					WHEN	239	=>	bit_input<='1';
					WHEN	240	=>	bit_input<='1';
					WHEN	241	=>	bit_input<='1';
					WHEN	242	=>	bit_input<='1';
					WHEN	243	=>	bit_input<='1';
					WHEN	244	=>	bit_input<='1';
					WHEN	245	=>	bit_input<='1';
					WHEN	246	=>	bit_input<='1';
					WHEN	247	=>	bit_input<='1';
					WHEN	248	=>	bit_input<='1';
					WHEN	249	=>	bit_input<='1';
					WHEN	250	=>	bit_input<='1';
					WHEN	251	=>	bit_input<='1';
					WHEN	252	=>	bit_input<='1';
					WHEN	253	=>	bit_input<='1';
					WHEN	254	=>	bit_input<='1';
					WHEN	255	=>	bit_input<='1';
					WHEN	256	=>	bit_input<='1';
					WHEN	257	=>	bit_input<='1';
					WHEN	258	=>	bit_input<='1';
					WHEN	259	=>	bit_input<='1';
					WHEN	260	=>	bit_input<='1';
					WHEN	261	=>	bit_input<='1';
					WHEN	262	=>	bit_input<='1';
					WHEN	263	=>	bit_input<='1';
					WHEN	264	=>	bit_input<='1';
					WHEN	265	=>	bit_input<='1';
					WHEN	266	=>	bit_input<='1';
					WHEN	267	=>	bit_input<='1';
					WHEN	268	=>	bit_input<='1';
					WHEN	269	=>	bit_input<='1';
					WHEN	270	=>	bit_input<='1';
					WHEN	271	=>	bit_input<='1';
					WHEN	272	=>	bit_input<='1';
					WHEN	273	=>	bit_input<='1';
					WHEN	274	=>	bit_input<='1';
					WHEN	275	=>	bit_input<='1';
					WHEN	276	=>	bit_input<='1';
					WHEN	277	=>	bit_input<='1';
					WHEN	278	=>	bit_input<='1';
					WHEN	279	=>	bit_input<='1';
					WHEN	280	=>	bit_input<='1';
					WHEN	281	=>	bit_input<='1';
					WHEN	282	=>	bit_input<='1';
					WHEN	283	=>	bit_input<='1';
					WHEN	284	=>	bit_input<='1';
					WHEN	285	=>	bit_input<='1';
					WHEN	286	=>	bit_input<='1';
					WHEN	287	=>	bit_input<='1';
					WHEN	288	=>	bit_input<='1';
					WHEN	289	=>	bit_input<='1';
					WHEN	290	=>	bit_input<='1';
					WHEN	291	=>	bit_input<='1';
					WHEN	292	=>	bit_input<='1';
					WHEN	293	=>	bit_input<='1';
					WHEN	294	=>	bit_input<='1';
					WHEN	295	=>	bit_input<='1';
					WHEN	296	=>	bit_input<='1';
					WHEN	297	=>	bit_input<='1';
					WHEN	298	=>	bit_input<='1';
					WHEN	299	=>	bit_input<='1';
					WHEN	300	=>	bit_input<='1';
					WHEN	301	=>	bit_input<='1';
					WHEN	302	=>	bit_input<='1';
					WHEN	303	=>	bit_input<='1';
					WHEN	304	=>	bit_input<='1';
					WHEN	305	=>	bit_input<='1';
					WHEN	306	=>	bit_input<='1';
					WHEN	307	=>	bit_input<='1';
					WHEN	308	=>	bit_input<='1';
					WHEN	309	=>	bit_input<='1';
					WHEN	310	=>	bit_input<='1';
					WHEN	311	=>	bit_input<='1';
					WHEN	312	=>	bit_input<='1';
					WHEN	313	=>	bit_input<='1';
					WHEN	314	=>	bit_input<='1';
					WHEN	315	=>	bit_input<='1';
					WHEN	316	=>	bit_input<='1';
					WHEN	317	=>	bit_input<='1';
					WHEN	318	=>	bit_input<='1';
					WHEN	319	=>	bit_input<='1';
					WHEN	320	=>	bit_input<='1';
					WHEN	321	=>	bit_input<='1';
					WHEN	322	=>	bit_input<='1';
					WHEN	323	=>	bit_input<='1';
					WHEN	324	=>	bit_input<='1';
					WHEN	325	=>	bit_input<='1';
					WHEN	326	=>	bit_input<='1';
					WHEN	327	=>	bit_input<='1';
					WHEN	328	=>	bit_input<='1';
					WHEN	329	=>	bit_input<='1';
					WHEN	330	=>	bit_input<='1';
					WHEN	331	=>	bit_input<='1';
					WHEN	332	=>	bit_input<='1';
					WHEN	333	=>	bit_input<='1';
					WHEN	334	=>	bit_input<='1';
					WHEN	335	=>	bit_input<='1';
					WHEN	336	=>	bit_input<='1';
					WHEN	337	=>	bit_input<='1';
					WHEN	338	=>	bit_input<='1';
					WHEN	339	=>	bit_input<='1';
					WHEN	340	=>	bit_input<='1';
					WHEN	341	=>	bit_input<='1';
					WHEN	342	=>	bit_input<='1';
					WHEN	343	=>	bit_input<='1';
					WHEN	344	=>	bit_input<='1';
					WHEN	345	=>	bit_input<='1';
					WHEN	346	=>	bit_input<='1';
					WHEN	347	=>	bit_input<='1';
					WHEN	348	=>	bit_input<='1';
					WHEN	349	=>	bit_input<='1';
					WHEN	350	=>	bit_input<='1';
					WHEN	351	=>	bit_input<='1';
					WHEN	352	=>	bit_input<='1';
					WHEN	353	=>	bit_input<='1';
					WHEN	354	=>	bit_input<='1';
					WHEN	355	=>	bit_input<='1';
					WHEN	356	=>	bit_input<='1';
					WHEN	357	=>	bit_input<='1';
					WHEN	358	=>	bit_input<='1';
					WHEN	359	=>	bit_input<='1';
					WHEN	360	=>	bit_input<='1';
					WHEN	361	=>	bit_input<='1';
					WHEN	362	=>	bit_input<='1';
					WHEN	363	=>	bit_input<='1';
					WHEN	364	=>	bit_input<='1';
					WHEN	365	=>	bit_input<='1';
					WHEN	366	=>	bit_input<='1';
					WHEN	367	=>	bit_input<='1';
					WHEN	368	=>	bit_input<='1';
					WHEN	369	=>	bit_input<='1';
					WHEN	370	=>	bit_input<='1';
					WHEN	371	=>	bit_input<='1';
					WHEN	372	=>	bit_input<='1';
					WHEN	373	=>	bit_input<='1';
					WHEN	374	=>	bit_input<='1';
					WHEN	375	=>	bit_input<='1';
					WHEN	376	=>	bit_input<='1';
					WHEN	377	=>	bit_input<='1';
					WHEN	378	=>	bit_input<='1';
					WHEN	379	=>	bit_input<='1';
					WHEN	380	=>	bit_input<='1';
					WHEN	381	=>	bit_input<='1';
					WHEN	382	=>	bit_input<='1';
					WHEN	383	=>	bit_input<='1';
					WHEN	384	=>	bit_input<='1';
					WHEN	385	=>	bit_input<='1';
					WHEN	386	=>	bit_input<='1';
					WHEN	387	=>	bit_input<='1';
					WHEN	388	=>	bit_input<='1';
					WHEN	389	=>	bit_input<='1';
					WHEN	390	=>	bit_input<='1';
					WHEN	391	=>	bit_input<='1';
					WHEN	392	=>	bit_input<='1';
					WHEN	393	=>	bit_input<='1';
					WHEN	394	=>	bit_input<='1';
					WHEN	395	=>	bit_input<='1';
					WHEN	396	=>	bit_input<='1';
					WHEN	397	=>	bit_input<='1';
					WHEN	398	=>	bit_input<='1';
					WHEN	399	=>	bit_input<='1';
					WHEN	400	=>	bit_input<='1';
					WHEN	401	=>	bit_input<='1';
					WHEN	402	=>	bit_input<='1';
					WHEN	403	=>	bit_input<='1';
					WHEN	404	=>	bit_input<='1';
					WHEN	405	=>	bit_input<='1';
					WHEN	406	=>	bit_input<='1';
					WHEN	407	=>	bit_input<='1';
					WHEN	408	=>	bit_input<='1';
					WHEN	409	=>	bit_input<='1';
					WHEN	410	=>	bit_input<='1';
					WHEN	411	=>	bit_input<='1';
					WHEN	412	=>	bit_input<='1';
					WHEN	413	=>	bit_input<='1';
					WHEN	414	=>	bit_input<='1';
					WHEN	415	=>	bit_input<='1';
					WHEN	416	=>	bit_input<='1';
					WHEN	417	=>	bit_input<='1';
					WHEN	418	=>	bit_input<='1';
					WHEN	419	=>	bit_input<='1';
					WHEN	420	=>	bit_input<='1';
					WHEN	421	=>	bit_input<='1';
					WHEN	422	=>	bit_input<='1';
					WHEN	423	=>	bit_input<='1';
					WHEN	424	=>	bit_input<='1';
					WHEN	425	=>	bit_input<='1';
					WHEN	426	=>	bit_input<='1';
					WHEN	427	=>	bit_input<='1';
					WHEN	428	=>	bit_input<='1';
					WHEN	429	=>	bit_input<='1';
					WHEN	430	=>	bit_input<='1';
					WHEN	431	=>	bit_input<='1';
					WHEN	432	=>	bit_input<='1';
					WHEN	433	=>	bit_input<='1';
					WHEN	434	=>	bit_input<='1';
					WHEN	435	=>	bit_input<='1';
					WHEN	436	=>	bit_input<='1';
					WHEN	437	=>	bit_input<='1';
					WHEN	438	=>	bit_input<='1';
					WHEN	439	=>	bit_input<='1';
					WHEN	440	=>	bit_input<='1';
					WHEN	441	=>	bit_input<='1';
					WHEN	442	=>	bit_input<='1';
					WHEN	443	=>	bit_input<='1';
					WHEN	444	=>	bit_input<='1';
					WHEN	445	=>	bit_input<='1';
					WHEN	446	=>	bit_input<='1';
					WHEN	447	=>	bit_input<='1';
					WHEN	448	=>	bit_input<='1';
					WHEN	449	=>	bit_input<='1';
					WHEN	450	=>	bit_input<='1';
					WHEN	451	=>	bit_input<='1';
					WHEN	452	=>	bit_input<='1';
					WHEN	453	=>	bit_input<='1';
					WHEN	454	=>	bit_input<='1';
					WHEN	455	=>	bit_input<='1';
					WHEN	456	=>	bit_input<='1';
					WHEN	457	=>	bit_input<='1';
					WHEN	458	=>	bit_input<='1';
					WHEN	459	=>	bit_input<='1';
					WHEN	460	=>	bit_input<='1';
					WHEN	461	=>	bit_input<='1';
					WHEN	462	=>	bit_input<='1';
					WHEN	463	=>	bit_input<='1';
					WHEN	464	=>	bit_input<='1';
					WHEN	465	=>	bit_input<='1';
					WHEN	466	=>	bit_input<='1';
					WHEN	467	=>	bit_input<='1';
					WHEN	468	=>	bit_input<='1';
					WHEN	469	=>	bit_input<='1';
					WHEN	470	=>	bit_input<='1';
					WHEN	471	=>	bit_input<='1';
					WHEN	472	=>	bit_input<='1';
					WHEN	473	=>	bit_input<='1';
					WHEN	474	=>	bit_input<='1';
					WHEN	475	=>	bit_input<='1';
					WHEN	476	=>	bit_input<='1';
					WHEN	477	=>	bit_input<='1';
					WHEN	478	=>	bit_input<='1';
					WHEN	479	=>	bit_input<='1';
					WHEN	480	=>	bit_input<='1';
					WHEN	481	=>	bit_input<='1';
					WHEN	482	=>	bit_input<='1';
					WHEN	483	=>	bit_input<='1';
					WHEN	484	=>	bit_input<='1';
					WHEN	485	=>	bit_input<='1';
					WHEN	486	=>	bit_input<='1';
					WHEN	487	=>	bit_input<='1';
					WHEN	488	=>	bit_input<='1';
					WHEN	489	=>	bit_input<='1';
					WHEN	490	=>	bit_input<='1';
					WHEN	491	=>	bit_input<='1';
					WHEN	492	=>	bit_input<='1';
					WHEN	493	=>	bit_input<='1';
					WHEN	494	=>	bit_input<='1';
					WHEN	495	=>	bit_input<='1';
					WHEN	496	=>	bit_input<='1';
					WHEN	497	=>	bit_input<='1';
					WHEN	498	=>	bit_input<='1';
					WHEN	499	=>	bit_input<='1';
					WHEN	500	=>	bit_input<='1';
					WHEN	501	=>	bit_input<='1';
					WHEN	502	=>	bit_input<='1';
					WHEN	503	=>	bit_input<='1';
					WHEN	504	=>	bit_input<='1';
					WHEN	505	=>	bit_input<='1';
					WHEN	506	=>	bit_input<='1';
					WHEN	507	=>	bit_input<='1';
					WHEN	508	=>	bit_input<='1';
					WHEN	509	=>	bit_input<='1';
					WHEN	510	=>	bit_input<='1';
					WHEN	511	=>	bit_input<='1';
					WHEN	512	=>	bit_input<='1';
					WHEN	513	=>	bit_input<='1';
					WHEN	514	=>	bit_input<='1';
					WHEN	515	=>	bit_input<='1';
					WHEN	516	=>	bit_input<='1';
					WHEN	517	=>	bit_input<='1';
					WHEN	518	=>	bit_input<='1';
					WHEN	519	=>	bit_input<='1';
					WHEN	520	=>	bit_input<='1';
					WHEN	521	=>	bit_input<='1';
					WHEN	522	=>	bit_input<='1';
					WHEN	523	=>	bit_input<='1';
					WHEN	524	=>	bit_input<='1';
					WHEN	525	=>	bit_input<='1';
					WHEN	526	=>	bit_input<='1';
					WHEN	527	=>	bit_input<='1';
					WHEN	528	=>	bit_input<='1';
					WHEN	529	=>	bit_input<='1';
					WHEN	530	=>	bit_input<='1';
					WHEN	531	=>	bit_input<='1';
					WHEN	532	=>	bit_input<='1';
					WHEN	533	=>	bit_input<='1';
					WHEN	534	=>	bit_input<='1';
					WHEN	535	=>	bit_input<='1';
					WHEN	536	=>	bit_input<='1';
					WHEN	537	=>	bit_input<='1';
					WHEN	538	=>	bit_input<='1';
					WHEN	539	=>	bit_input<='1';
					WHEN	540	=>	bit_input<='1';
					WHEN	541	=>	bit_input<='1';
					WHEN	542	=>	bit_input<='1';
					WHEN	543	=>	bit_input<='1';
					WHEN	544	=>	bit_input<='1';
					WHEN	545	=>	bit_input<='1';
					WHEN	546	=>	bit_input<='1';
					WHEN	547	=>	bit_input<='1';
					WHEN	548	=>	bit_input<='1';
					WHEN	549	=>	bit_input<='1';
					WHEN	550	=>	bit_input<='1';
					WHEN	551	=>	bit_input<='1';
					WHEN	552	=>	bit_input<='1';
					WHEN	553	=>	bit_input<='1';
					WHEN	554	=>	bit_input<='1';
					WHEN	555	=>	bit_input<='1';
					WHEN	556	=>	bit_input<='1';
					WHEN	557	=>	bit_input<='1';
					WHEN	558	=>	bit_input<='1';
					WHEN	559	=>	bit_input<='1';
					WHEN	560	=>	bit_input<='1';
					WHEN	561	=>	bit_input<='1';
					WHEN	562	=>	bit_input<='1';
					WHEN	563	=>	bit_input<='1';
					WHEN	564	=>	bit_input<='1';
					WHEN	565	=>	bit_input<='1';
					WHEN	566	=>	bit_input<='1';
					WHEN	567	=>	bit_input<='1';
					WHEN	568	=>	bit_input<='1';
					WHEN	569	=>	bit_input<='1';
					WHEN	570	=>	bit_input<='1';
					WHEN	571	=>	bit_input<='1';
					WHEN	572	=>	bit_input<='1';
					WHEN	573	=>	bit_input<='1';
					WHEN	574	=>	bit_input<='1';
					WHEN	575	=>	bit_input<='1';
					WHEN	576	=>	bit_input<='1';
					WHEN	577	=>	bit_input<='1';
					WHEN	578	=>	bit_input<='1';
					WHEN	579	=>	bit_input<='1';
					WHEN	580	=>	bit_input<='1';
					WHEN	581	=>	bit_input<='1';
					WHEN	582	=>	bit_input<='1';
					WHEN	583	=>	bit_input<='1';
					WHEN	584	=>	bit_input<='1';
					WHEN	585	=>	bit_input<='1';
					WHEN	586	=>	bit_input<='1';
					WHEN	587	=>	bit_input<='1';
					WHEN	588	=>	bit_input<='1';
					WHEN	589	=>	bit_input<='1';
					WHEN	590	=>	bit_input<='1';
					WHEN	591	=>	bit_input<='1';
					WHEN	592	=>	bit_input<='1';
					WHEN	593	=>	bit_input<='1';
					WHEN	594	=>	bit_input<='1';
					WHEN	595	=>	bit_input<='1';
					WHEN	596	=>	bit_input<='1';
					WHEN	597	=>	bit_input<='1';
					WHEN	598	=>	bit_input<='1';
					WHEN	599	=>	bit_input<='1';
					WHEN	600	=>	bit_input<='1';
					WHEN	601	=>	bit_input<='1';
					WHEN	602	=>	bit_input<='1';
					WHEN	603	=>	bit_input<='1';
					WHEN	604	=>	bit_input<='1';
					WHEN	605	=>	bit_input<='1';
					WHEN	606	=>	bit_input<='1';
					WHEN	607	=>	bit_input<='1';
					WHEN	608	=>	bit_input<='1';
					WHEN	609	=>	bit_input<='1';
					WHEN	610	=>	bit_input<='1';
					WHEN	611	=>	bit_input<='1';
					WHEN	612	=>	bit_input<='1';
					WHEN	613	=>	bit_input<='1';
					WHEN	614	=>	bit_input<='1';
					WHEN	615	=>	bit_input<='1';
					WHEN	616	=>	bit_input<='1';
					WHEN	617	=>	bit_input<='1';
					WHEN	618	=>	bit_input<='1';
					WHEN	619	=>	bit_input<='1';
					WHEN	620	=>	bit_input<='1';
					WHEN	621	=>	bit_input<='1';
					WHEN	622	=>	bit_input<='1';
					WHEN	623	=>	bit_input<='1';
					WHEN	624	=>	bit_input<='1';
					WHEN	625	=>	bit_input<='1';
					WHEN	626	=>	bit_input<='1';
					WHEN	627	=>	bit_input<='1';
					WHEN	628	=>	bit_input<='1';
					WHEN	629	=>	bit_input<='1';
					WHEN	630	=>	bit_input<='1';
					WHEN	631	=>	bit_input<='1';
					WHEN	632	=>	bit_input<='1';
					WHEN	633	=>	bit_input<='1';
					WHEN	634	=>	bit_input<='1';
					WHEN	635	=>	bit_input<='1';
					WHEN	636	=>	bit_input<='1';
					WHEN	637	=>	bit_input<='1';
					WHEN	638	=>	bit_input<='1';
					WHEN	639	=>	bit_input<='1';
					WHEN	640	=>	bit_input<='1';
					WHEN	641	=>	bit_input<='1';
					WHEN	642	=>	bit_input<='1';
					WHEN	643	=>	bit_input<='1';
					WHEN	644	=>	bit_input<='1';
					WHEN	645	=>	bit_input<='1';
					WHEN	646	=>	bit_input<='1';
					WHEN	647	=>	bit_input<='1';
					WHEN	648	=>	bit_input<='1';
					WHEN	649	=>	bit_input<='1';
					WHEN	650	=>	bit_input<='1';
					WHEN	651	=>	bit_input<='1';
					WHEN	652	=>	bit_input<='1';
					WHEN	653	=>	bit_input<='1';
					WHEN	654	=>	bit_input<='1';
					WHEN	655	=>	bit_input<='1';
					WHEN	656	=>	bit_input<='1';
					WHEN	657	=>	bit_input<='1';
					WHEN	658	=>	bit_input<='1';
					WHEN	659	=>	bit_input<='1';
					WHEN	660	=>	bit_input<='1';
					WHEN	661	=>	bit_input<='1';
					WHEN	662	=>	bit_input<='1';
					WHEN	663	=>	bit_input<='1';
					WHEN	664	=>	bit_input<='1';
					WHEN	665	=>	bit_input<='1';
					WHEN	666	=>	bit_input<='1';
					WHEN	667	=>	bit_input<='1';
					WHEN	668	=>	bit_input<='1';
					WHEN	669	=>	bit_input<='1';
					WHEN	670	=>	bit_input<='1';
					WHEN	671	=>	bit_input<='1';
					WHEN	672	=>	bit_input<='1';
					WHEN	673	=>	bit_input<='1';
					WHEN	674	=>	bit_input<='1';
					WHEN	675	=>	bit_input<='1';
					WHEN	676	=>	bit_input<='1';
					WHEN	677	=>	bit_input<='1';
					WHEN	678	=>	bit_input<='1';
					WHEN	679	=>	bit_input<='1';
					WHEN	680	=>	bit_input<='1';
					WHEN	681	=>	bit_input<='1';
					WHEN	682	=>	bit_input<='1';
					WHEN	683	=>	bit_input<='1';
					WHEN	684	=>	bit_input<='1';
					WHEN	685	=>	bit_input<='1';
					WHEN	686	=>	bit_input<='1';
					WHEN	687	=>	bit_input<='1';
					WHEN	688	=>	bit_input<='1';
					WHEN	689	=>	bit_input<='1';
					WHEN	690	=>	bit_input<='1';
					WHEN	691	=>	bit_input<='1';
					WHEN	692	=>	bit_input<='1';
					WHEN	693	=>	bit_input<='1';
					WHEN	694	=>	bit_input<='1';
					WHEN	695	=>	bit_input<='1';
					WHEN	696	=>	bit_input<='1';
					WHEN	697	=>	bit_input<='1';
					WHEN	698	=>	bit_input<='1';
					WHEN	699	=>	bit_input<='1';
					WHEN	700	=>	bit_input<='1';
					WHEN	701	=>	bit_input<='1';
					WHEN	702	=>	bit_input<='1';
					WHEN	703	=>	bit_input<='1';
					WHEN	704	=>	bit_input<='1';
					WHEN	705	=>	bit_input<='1';
					WHEN	706	=>	bit_input<='1';
					WHEN	707	=>	bit_input<='1';
					WHEN	708	=>	bit_input<='1';
					WHEN	709	=>	bit_input<='1';
					WHEN	710	=>	bit_input<='1';
					WHEN	711	=>	bit_input<='1';
					WHEN	712	=>	bit_input<='1';
					WHEN	713	=>	bit_input<='1';
					WHEN	714	=>	bit_input<='1';
					WHEN	715	=>	bit_input<='1';
					WHEN	716	=>	bit_input<='1';
					WHEN	717	=>	bit_input<='1';
					WHEN	718	=>	bit_input<='1';
					WHEN	719	=>	bit_input<='1';
					WHEN	720	=>	bit_input<='1';
					WHEN	721	=>	bit_input<='1';
					WHEN	722	=>	bit_input<='1';
					WHEN	723	=>	bit_input<='1';
					WHEN	724	=>	bit_input<='1';
					WHEN	725	=>	bit_input<='1';
					WHEN	726	=>	bit_input<='1';
					WHEN	727	=>	bit_input<='1';
					WHEN	728	=>	bit_input<='1';
					WHEN	729	=>	bit_input<='1';
					WHEN	730	=>	bit_input<='1';
					WHEN	731	=>	bit_input<='1';
					WHEN	732	=>	bit_input<='1';
					WHEN	733	=>	bit_input<='1';
					WHEN	734	=>	bit_input<='1';
					WHEN	735	=>	bit_input<='1';
					WHEN	736	=>	bit_input<='1';
					WHEN	737	=>	bit_input<='1';
					WHEN	738	=>	bit_input<='1';
					WHEN	739	=>	bit_input<='1';
					WHEN	740	=>	bit_input<='1';
					WHEN	741	=>	bit_input<='1';
					WHEN	742	=>	bit_input<='1';
					WHEN	743	=>	bit_input<='1';
					WHEN	744	=>	bit_input<='1';
					WHEN	745	=>	bit_input<='1';
					WHEN	746	=>	bit_input<='1';
					WHEN	747	=>	bit_input<='1';
					WHEN	748	=>	bit_input<='1';
					WHEN	749	=>	bit_input<='1';
					WHEN	750	=>	bit_input<='1';
					WHEN	751	=>	bit_input<='1';
					WHEN	752	=>	bit_input<='1';
					WHEN	753	=>	bit_input<='1';
					WHEN	754	=>	bit_input<='1';
					WHEN	755	=>	bit_input<='1';
					WHEN	756	=>	bit_input<='1';
					WHEN	757	=>	bit_input<='1';
					WHEN	758	=>	bit_input<='1';
					WHEN	759	=>	bit_input<='1';
					WHEN	760	=>	bit_input<='1';
					WHEN	761	=>	bit_input<='1';
					WHEN	762	=>	bit_input<='1';
					WHEN	763	=>	bit_input<='1';
					WHEN	764	=>	bit_input<='1';
					WHEN	765	=>	bit_input<='1';
					WHEN	766	=>	bit_input<='1';
					WHEN	767	=>	bit_input<='1';
					WHEN	768	=>	bit_input<='1';
					WHEN	769	=>	bit_input<='1';
					WHEN	770	=>	bit_input<='1';
					WHEN	771	=>	bit_input<='1';
					WHEN	772	=>	bit_input<='1';
					WHEN	773	=>	bit_input<='1';
					WHEN	774	=>	bit_input<='1';
					WHEN	775	=>	bit_input<='1';
					WHEN	776	=>	bit_input<='1';
					WHEN	777	=>	bit_input<='1';
					WHEN	778	=>	bit_input<='1';
					WHEN	779	=>	bit_input<='1';
					WHEN	780	=>	bit_input<='1';
					WHEN	781	=>	bit_input<='1';
					WHEN	782	=>	bit_input<='1';
					WHEN	783	=>	bit_input<='1';
					WHEN	784	=>	bit_input<='1';
					WHEN	785	=>	bit_input<='1';
					WHEN	786	=>	bit_input<='1';
					WHEN	787	=>	bit_input<='1';
					WHEN	788	=>	bit_input<='1';
					WHEN	789	=>	bit_input<='1';
					WHEN	790	=>	bit_input<='1';
					WHEN	791	=>	bit_input<='1';
					WHEN	792	=>	bit_input<='1';
					WHEN	793	=>	bit_input<='1';
					WHEN	794	=>	bit_input<='1';
					WHEN	795	=>	bit_input<='1';
					WHEN	796	=>	bit_input<='1';
					WHEN	797	=>	bit_input<='1';
					WHEN	798	=>	bit_input<='1';
					WHEN	799	=>	bit_input<='1';
					WHEN	800	=>	bit_input<='1';
					WHEN	801	=>	bit_input<='1';
					WHEN	802	=>	bit_input<='1';
					WHEN	803	=>	bit_input<='1';
					WHEN	804	=>	bit_input<='1';
					WHEN	805	=>	bit_input<='1';
					WHEN	806	=>	bit_input<='1';
					WHEN	807	=>	bit_input<='1';
					WHEN	808	=>	bit_input<='1';
					WHEN	809	=>	bit_input<='1';
					WHEN	810	=>	bit_input<='1';
					WHEN	811	=>	bit_input<='1';
					WHEN	812	=>	bit_input<='1';
					WHEN	813	=>	bit_input<='1';
					WHEN	814	=>	bit_input<='1';
					WHEN	815	=>	bit_input<='1';
					WHEN	816	=>	bit_input<='1';
					WHEN	817	=>	bit_input<='1';
					WHEN	818	=>	bit_input<='1';
					WHEN	819	=>	bit_input<='1';
					WHEN	820	=>	bit_input<='1';
					WHEN	821	=>	bit_input<='1';
					WHEN	822	=>	bit_input<='1';
					WHEN	823	=>	bit_input<='1';
					WHEN	824	=>	bit_input<='1';
					WHEN	825	=>	bit_input<='1';
					WHEN	826	=>	bit_input<='1';
					WHEN	827	=>	bit_input<='1';
					WHEN	828	=>	bit_input<='1';
					WHEN	829	=>	bit_input<='1';
					WHEN	830	=>	bit_input<='1';
					WHEN	831	=>	bit_input<='1';
					WHEN	832	=>	bit_input<='1';
					WHEN	833	=>	bit_input<='1';
					WHEN	834	=>	bit_input<='1';
					WHEN	835	=>	bit_input<='1';
					WHEN	836	=>	bit_input<='1';
					WHEN	837	=>	bit_input<='1';
					WHEN	838	=>	bit_input<='1';
					WHEN	839	=>	bit_input<='1';
					WHEN	840	=>	bit_input<='1';
					WHEN	841	=>	bit_input<='1';
					WHEN	842	=>	bit_input<='1';
					WHEN	843	=>	bit_input<='1';
					WHEN	844	=>	bit_input<='1';
					WHEN	845	=>	bit_input<='1';
					WHEN	846	=>	bit_input<='1';
					WHEN	847	=>	bit_input<='1';
					WHEN	848	=>	bit_input<='1';
					WHEN	849	=>	bit_input<='1';
					WHEN	850	=>	bit_input<='1';
					WHEN	851	=>	bit_input<='1';
					WHEN	852	=>	bit_input<='1';
					WHEN	853	=>	bit_input<='1';
					WHEN	854	=>	bit_input<='1';
					WHEN	855	=>	bit_input<='1';
					WHEN	856	=>	bit_input<='1';
					WHEN	857	=>	bit_input<='1';
					WHEN	858	=>	bit_input<='1';
					WHEN	859	=>	bit_input<='1';
					WHEN	860	=>	bit_input<='1';
					WHEN	861	=>	bit_input<='1';
					WHEN	862	=>	bit_input<='1';
					WHEN	863	=>	bit_input<='1';
					WHEN	864	=>	bit_input<='1';
					WHEN	865	=>	bit_input<='1';
					WHEN	866	=>	bit_input<='1';
					WHEN	867	=>	bit_input<='1';
					WHEN	868	=>	bit_input<='1';
					WHEN	869	=>	bit_input<='1';
					WHEN	870	=>	bit_input<='1';
					WHEN	871	=>	bit_input<='1';
					WHEN	872	=>	bit_input<='1';
					WHEN	873	=>	bit_input<='1';
					WHEN	874	=>	bit_input<='1';
					WHEN	875	=>	bit_input<='1';
					WHEN	876	=>	bit_input<='1';
					WHEN	877	=>	bit_input<='1';
					WHEN	878	=>	bit_input<='1';
					WHEN	879	=>	bit_input<='1';
					WHEN	880	=>	bit_input<='1';
					WHEN	881	=>	bit_input<='1';
					WHEN	882	=>	bit_input<='1';
					WHEN	883	=>	bit_input<='1';
					WHEN	884	=>	bit_input<='1';
					WHEN	885	=>	bit_input<='1';
					WHEN	886	=>	bit_input<='1';
					WHEN	887	=>	bit_input<='1';
					WHEN	888	=>	bit_input<='1';
					WHEN	889	=>	bit_input<='1';
					WHEN	890	=>	bit_input<='1';
					WHEN	891	=>	bit_input<='1';
					WHEN	892	=>	bit_input<='1';
					WHEN	893	=>	bit_input<='1';
					WHEN	894	=>	bit_input<='1';
					WHEN	895	=>	bit_input<='1';
					WHEN	896	=>	bit_input<='1';
					WHEN	897	=>	bit_input<='1';
					WHEN	898	=>	bit_input<='1';
					WHEN	899	=>	bit_input<='1';
					WHEN	900	=>	bit_input<='1';
					WHEN	901	=>	bit_input<='1';
					WHEN	902	=>	bit_input<='1';
					WHEN	903	=>	bit_input<='1';
					WHEN	904	=>	bit_input<='1';
					WHEN	905	=>	bit_input<='1';
					WHEN	906	=>	bit_input<='1';
					WHEN	907	=>	bit_input<='1';
					WHEN	908	=>	bit_input<='1';
					WHEN	909	=>	bit_input<='1';
					WHEN	910	=>	bit_input<='1';
					WHEN	911	=>	bit_input<='1';
					WHEN	912	=>	bit_input<='1';
					WHEN	913	=>	bit_input<='1';
					WHEN	914	=>	bit_input<='1';
					WHEN	915	=>	bit_input<='1';
					WHEN	916	=>	bit_input<='1';
					WHEN	917	=>	bit_input<='1';
					WHEN	918	=>	bit_input<='1';
					WHEN	919	=>	bit_input<='1';
					WHEN	920	=>	bit_input<='1';
					WHEN	921	=>	bit_input<='1';
					WHEN	922	=>	bit_input<='1';
					WHEN	923	=>	bit_input<='1';
					WHEN	924	=>	bit_input<='1';
					WHEN	925	=>	bit_input<='1';
					WHEN	926	=>	bit_input<='1';
					WHEN	927	=>	bit_input<='1';
					WHEN	928	=>	bit_input<='1';
					WHEN	929	=>	bit_input<='1';
					WHEN	930	=>	bit_input<='1';
					WHEN	931	=>	bit_input<='1';
					WHEN	932	=>	bit_input<='1';
					WHEN	933	=>	bit_input<='1';
					WHEN	934	=>	bit_input<='1';
					WHEN	935	=>	bit_input<='1';
					WHEN	936	=>	bit_input<='1';
					WHEN	937	=>	bit_input<='1';
					WHEN	938	=>	bit_input<='1';
					WHEN	939	=>	bit_input<='1';
					WHEN	940	=>	bit_input<='1';
					WHEN	941	=>	bit_input<='1';
					WHEN	942	=>	bit_input<='1';
					WHEN	943	=>	bit_input<='1';
					WHEN	944	=>	bit_input<='1';
					WHEN	945	=>	bit_input<='1';
					WHEN	946	=>	bit_input<='1';
					WHEN	947	=>	bit_input<='1';
					WHEN	948	=>	bit_input<='1';
					WHEN	949	=>	bit_input<='1';
					WHEN	950	=>	bit_input<='1';
					WHEN	951	=>	bit_input<='1';
					WHEN	952	=>	bit_input<='1';
					WHEN	953	=>	bit_input<='1';
					WHEN	954	=>	bit_input<='1';
					WHEN	955	=>	bit_input<='1';
					WHEN	956	=>	bit_input<='1';
					WHEN	957	=>	bit_input<='1';
					WHEN	958	=>	bit_input<='1';
					WHEN	959	=>	bit_input<='1';
					WHEN	960	=>	bit_input<='1';
					WHEN	961	=>	bit_input<='1';
					WHEN	962	=>	bit_input<='1';
					WHEN	963	=>	bit_input<='1';
					WHEN	964	=>	bit_input<='1';
					WHEN	965	=>	bit_input<='1';
					WHEN	966	=>	bit_input<='1';
					WHEN	967	=>	bit_input<='1';
					WHEN	968	=>	bit_input<='1';
					WHEN	969	=>	bit_input<='1';
					WHEN	970	=>	bit_input<='1';
					WHEN	971	=>	bit_input<='1';
					WHEN	972	=>	bit_input<='1';
					WHEN	973	=>	bit_input<='1';
					WHEN	974	=>	bit_input<='1';
					WHEN	975	=>	bit_input<='1';
					WHEN	976	=>	bit_input<='1';
					WHEN	977	=>	bit_input<='1';
					WHEN	978	=>	bit_input<='1';
					WHEN	979	=>	bit_input<='1';
					WHEN	980	=>	bit_input<='1';
					WHEN	981	=>	bit_input<='1';
					WHEN	982	=>	bit_input<='1';
					WHEN	983	=>	bit_input<='1';
					WHEN	984	=>	bit_input<='1';
					WHEN	985	=>	bit_input<='1';
					WHEN	986	=>	bit_input<='1';
					WHEN	987	=>	bit_input<='1';
					WHEN	988	=>	bit_input<='1';
					WHEN	989	=>	bit_input<='1';
					WHEN	990	=>	bit_input<='1';
					WHEN	991	=>	bit_input<='1';
					WHEN	992	=>	bit_input<='1';
					WHEN	993	=>	bit_input<='1';
					WHEN	994	=>	bit_input<='1';
					WHEN	995	=>	bit_input<='1';
					WHEN	996	=>	bit_input<='1';
					WHEN	997	=>	bit_input<='1';
					WHEN	998	=>	bit_input<='1';
					WHEN	999	=>	bit_input<='1';
					WHEN	1000	=>	bit_input<='1';
					WHEN	1001	=>	bit_input<='1';
					WHEN	1002	=>	bit_input<='1';
					WHEN	1003	=>	bit_input<='1';
					WHEN	1004	=>	bit_input<='1';
					WHEN	1005	=>	bit_input<='1';
					WHEN	1006	=>	bit_input<='1';
					WHEN	1007	=>	bit_input<='1';
					WHEN	1008	=>	bit_input<='1';
					WHEN	1009	=>	bit_input<='1';
					WHEN	1010	=>	bit_input<='1';
					WHEN	1011	=>	bit_input<='1';
					WHEN	1012	=>	bit_input<='1';
					WHEN	1013	=>	bit_input<='1';
					WHEN	1014	=>	bit_input<='1';
					WHEN	1015	=>	bit_input<='1';
					WHEN	1016	=>	bit_input<='1';
					WHEN	1017	=>	bit_input<='1';
					WHEN	1018	=>	bit_input<='1';
					WHEN	1019	=>	bit_input<='1';
					WHEN	1020	=>	bit_input<='1';
					WHEN	1021	=>	bit_input<='1';
					WHEN	1022	=>	bit_input<='1';
					WHEN	1023	=>	bit_input<='1';
					WHEN	1024	=>	bit_input<='1';

					-- starting output

					WHEN	1025	=>	bit_input<='Z';
					WHEN	1026	=>	bit_input<='Z';
					WHEN	1027	=>	bit_input<='Z';
					WHEN	1028	=>	bit_input<='Z';
					WHEN	1029	=>	bit_input<='Z';
					WHEN	1030	=>	bit_input<='Z';
					WHEN	1031	=>	bit_input<='Z';
					WHEN	1032	=>	bit_input<='Z';
					WHEN	1033	=>	bit_input<='Z';
					WHEN	1034	=>	bit_input<='Z';
					WHEN	1035	=>	bit_input<='Z';
					WHEN	1036	=>	bit_input<='Z';
					WHEN	1037	=>	bit_input<='Z';
					WHEN	1038	=>	bit_input<='Z';
					WHEN	1039	=>	bit_input<='Z';
					WHEN	1040	=>	bit_input<='Z';
					WHEN	1041	=>	bit_input<='Z';
					WHEN	1042	=>	bit_input<='Z';
					WHEN	1043	=>	bit_input<='Z';
					WHEN	1044	=>	bit_input<='Z';
					WHEN	1045	=>	bit_input<='Z';
					WHEN	1046	=>	bit_input<='Z';
					WHEN	1047	=>	bit_input<='Z';
					WHEN	1048	=>	bit_input<='Z';
					WHEN	1049	=>	bit_input<='Z';
					WHEN	1050	=>	bit_input<='Z';
					WHEN	1051	=>	bit_input<='Z';
					WHEN	1052	=>	bit_input<='Z';
					WHEN	1053	=>	bit_input<='Z';
					WHEN	1054	=>	bit_input<='Z';
					WHEN	1055	=>	bit_input<='Z';
					WHEN	1056	=>	bit_input<='Z';
					WHEN	1057	=>	bit_input<='Z';
					WHEN	1058	=>	bit_input<='Z';
					WHEN	1059	=>	bit_input<='Z';
					WHEN	1060	=>	bit_input<='Z';
					WHEN	1061	=>	bit_input<='Z';
					WHEN	1062	=>	bit_input<='Z';
					WHEN	1063	=>	bit_input<='Z';
					WHEN	1064	=>	bit_input<='Z';
					WHEN	1065	=>	bit_input<='Z';
					WHEN	1066	=>	bit_input<='Z';
					WHEN	1067	=>	bit_input<='Z';
					WHEN	1068	=>	bit_input<='Z';
					WHEN	1069	=>	bit_input<='Z';
					WHEN	1070	=>	bit_input<='Z';
					WHEN	1071	=>	bit_input<='Z';
					WHEN	1072	=>	bit_input<='Z';
					WHEN	1073	=>	bit_input<='Z';
					WHEN	1074	=>	bit_input<='Z';
					WHEN	1075	=>	bit_input<='Z';
					WHEN	1076	=>	bit_input<='Z';
					WHEN	1077	=>	bit_input<='Z';
					WHEN	1078	=>	bit_input<='Z';
					WHEN	1079	=>	bit_input<='Z';
					WHEN	1080	=>	bit_input<='Z';
					WHEN	1081	=>	bit_input<='Z';
					WHEN	1082	=>	bit_input<='Z';
					WHEN	1083	=>	bit_input<='Z';
					WHEN	1084	=>	bit_input<='Z';
					WHEN	1085	=>	bit_input<='Z';
					WHEN	1086	=>	bit_input<='Z';
					WHEN	1087	=>	bit_input<='Z';
					WHEN	1088	=>	bit_input<='Z';
					WHEN	1089	=>	bit_input<='Z';
					WHEN	1090	=>	bit_input<='Z';
					WHEN	1091	=>	bit_input<='Z';
					WHEN	1092	=>	bit_input<='Z';
					WHEN	1093	=>	bit_input<='Z';
					WHEN	1094	=>	bit_input<='Z';
					WHEN	1095	=>	bit_input<='Z';
					WHEN	1096	=>	bit_input<='Z';
					WHEN	1097	=>	bit_input<='Z';
					WHEN	1098	=>	bit_input<='Z';
					WHEN	1099	=>	bit_input<='Z';
					WHEN	1100	=>	bit_input<='Z';
					WHEN	1101	=>	bit_input<='Z';
					WHEN	1102	=>	bit_input<='Z';
					WHEN	1103	=>	bit_input<='Z';
					WHEN	1104	=>	bit_input<='Z';
					WHEN	1105	=>	bit_input<='Z';
					WHEN	1106	=>	bit_input<='Z';
					WHEN	1107	=>	bit_input<='Z';
					WHEN	1108	=>	bit_input<='Z';
					WHEN	1109	=>	bit_input<='Z';
					WHEN	1110	=>	bit_input<='Z';
					WHEN	1111	=>	bit_input<='Z';
					WHEN	1112	=>	bit_input<='Z';
					WHEN	1113	=>	bit_input<='Z';
					WHEN	1114	=>	bit_input<='Z';
					WHEN	1115	=>	bit_input<='Z';
					WHEN	1116	=>	bit_input<='Z';
					WHEN	1117	=>	bit_input<='Z';
					WHEN	1118	=>	bit_input<='Z';
					WHEN	1119	=>	bit_input<='Z';
					WHEN	1120	=>	bit_input<='Z';
					WHEN	1121	=>	bit_input<='Z';
					WHEN	1122	=>	bit_input<='Z';
					WHEN	1123	=>	bit_input<='Z';
					WHEN	1124	=>	bit_input<='Z';
					WHEN	1125	=>	bit_input<='Z';
					WHEN	1126	=>	bit_input<='Z';
					WHEN	1127	=>	bit_input<='Z';
					WHEN	1128	=>	bit_input<='Z';
					WHEN	1129	=>	bit_input<='Z';
					WHEN	1130	=>	bit_input<='Z';
					WHEN	1131	=>	bit_input<='Z';
					WHEN	1132	=>	bit_input<='Z';
					WHEN	1133	=>	bit_input<='Z';
					WHEN	1134	=>	bit_input<='Z';
					WHEN	1135	=>	bit_input<='Z';
					WHEN	1136	=>	bit_input<='Z';
					WHEN	1137	=>	bit_input<='Z';
					WHEN	1138	=>	bit_input<='Z';
					WHEN	1139	=>	bit_input<='Z';
					WHEN	1140	=>	bit_input<='Z';
					WHEN	1141	=>	bit_input<='Z';
					WHEN	1142	=>	bit_input<='Z';
					WHEN	1143	=>	bit_input<='Z';
					WHEN	1144	=>	bit_input<='Z';
					WHEN	1145	=>	bit_input<='Z';
					WHEN	1146	=>	bit_input<='Z';
					WHEN	1147	=>	bit_input<='Z';
					WHEN	1148	=>	bit_input<='Z';
					WHEN	1149	=>	bit_input<='Z';
					WHEN	1150	=>	bit_input<='Z';
					WHEN	1151	=>	bit_input<='Z';
					WHEN	1152	=>	bit_input<='Z';
					WHEN	1153	=>	bit_input<='Z';
					WHEN	1154	=>	bit_input<='Z';
					WHEN	1155	=>	bit_input<='Z';
					WHEN	1156	=>	bit_input<='Z';
					WHEN	1157	=>	bit_input<='Z';
					WHEN	1158	=>	bit_input<='Z';
					WHEN	1159	=>	bit_input<='Z';
					WHEN	1160	=>	bit_input<='Z';
					WHEN	1161	=>	bit_input<='Z';
					WHEN	1162	=>	bit_input<='Z';
					WHEN	1163	=>	bit_input<='Z';
					WHEN	1164	=>	bit_input<='Z';
					WHEN	1165	=>	bit_input<='Z';
					WHEN	1166	=>	bit_input<='Z';
					WHEN	1167	=>	bit_input<='Z';
					WHEN	1168	=>	bit_input<='Z';
					WHEN	1169	=>	bit_input<='Z';
					WHEN	1170	=>	bit_input<='Z';
					WHEN	1171	=>	bit_input<='Z';
					WHEN	1172	=>	bit_input<='Z';
					WHEN	1173	=>	bit_input<='Z';
					WHEN	1174	=>	bit_input<='Z';
					WHEN	1175	=>	bit_input<='Z';
					WHEN	1176	=>	bit_input<='Z';
					WHEN	1177	=>	bit_input<='Z';
					WHEN	1178	=>	bit_input<='Z';
					WHEN	1179	=>	bit_input<='Z';
					WHEN	1180	=>	bit_input<='Z';
					WHEN	1181	=>	bit_input<='Z';
					WHEN	1182	=>	bit_input<='Z';
					WHEN	1183	=>	bit_input<='Z';
					WHEN	1184	=>	bit_input<='Z';
					WHEN	1185	=>	bit_input<='Z';
					WHEN	1186	=>	bit_input<='Z';
					WHEN	1187	=>	bit_input<='Z';
					WHEN	1188	=>	bit_input<='Z';
					WHEN	1189	=>	bit_input<='Z';
					WHEN	1190	=>	bit_input<='Z';
					WHEN	1191	=>	bit_input<='Z';
					WHEN	1192	=>	bit_input<='Z';
					WHEN	1193	=>	bit_input<='Z';
					WHEN	1194	=>	bit_input<='Z';
					WHEN	1195	=>	bit_input<='Z';
					WHEN	1196	=>	bit_input<='Z';
					WHEN	1197	=>	bit_input<='Z';
					WHEN	1198	=>	bit_input<='Z';
					WHEN	1199	=>	bit_input<='Z';
					WHEN	1200	=>	bit_input<='Z';
					WHEN	1201	=>	bit_input<='Z';
					WHEN	1202	=>	bit_input<='Z';
					WHEN	1203	=>	bit_input<='Z';
					WHEN	1204	=>	bit_input<='Z';
					WHEN	1205	=>	bit_input<='Z';
					WHEN	1206	=>	bit_input<='Z';
					WHEN	1207	=>	bit_input<='Z';
					WHEN	1208	=>	bit_input<='Z';
					WHEN	1209	=>	bit_input<='Z';
					WHEN	1210	=>	bit_input<='Z';
					WHEN	1211	=>	bit_input<='Z';
					WHEN	1212	=>	bit_input<='Z';
					WHEN	1213	=>	bit_input<='Z';
					WHEN	1214	=>	bit_input<='Z';
					WHEN	1215	=>	bit_input<='Z';
					WHEN	1216	=>	bit_input<='Z';
					WHEN	1217	=>	bit_input<='Z';
					WHEN	1218	=>	bit_input<='Z';
					WHEN	1219	=>	bit_input<='Z';
					WHEN	1220	=>	bit_input<='Z';
					WHEN	1221	=>	bit_input<='Z';
					WHEN	1222	=>	bit_input<='Z';
					WHEN	1223	=>	bit_input<='Z';
					WHEN	1224	=>	bit_input<='Z';
					WHEN	1225	=>	bit_input<='Z';
					WHEN	1226	=>	bit_input<='Z';
					WHEN	1227	=>	bit_input<='Z';
					WHEN	1228	=>	bit_input<='Z';
					WHEN	1229	=>	bit_input<='Z';
					WHEN	1230	=>	bit_input<='Z';
					WHEN	1231	=>	bit_input<='Z';
					WHEN	1232	=>	bit_input<='Z';
					WHEN	1233	=>	bit_input<='Z';
					WHEN	1234	=>	bit_input<='Z';
					WHEN	1235	=>	bit_input<='Z';
					WHEN	1236	=>	bit_input<='Z';
					WHEN	1237	=>	bit_input<='Z';
					WHEN	1238	=>	bit_input<='Z';
					WHEN	1239	=>	bit_input<='Z';
					WHEN	1240	=>	bit_input<='Z';
					WHEN	1241	=>	bit_input<='Z';
					WHEN	1242	=>	bit_input<='Z';
					WHEN	1243	=>	bit_input<='Z';
					WHEN	1244	=>	bit_input<='Z';
					WHEN	1245	=>	bit_input<='Z';
					WHEN	1246	=>	bit_input<='Z';
					WHEN	1247	=>	bit_input<='Z';
					WHEN	1248	=>	bit_input<='Z';
					WHEN	1249	=>	bit_input<='Z';
					WHEN	1250	=>	bit_input<='Z';
					WHEN	1251	=>	bit_input<='Z';
					WHEN	1252	=>	bit_input<='Z';
					WHEN	1253	=>	bit_input<='Z';
					WHEN	1254	=>	bit_input<='Z';
					WHEN	1255	=>	bit_input<='Z';
					WHEN	1256	=>	bit_input<='Z';
					WHEN	1257	=>	bit_input<='Z';
					WHEN	1258	=>	bit_input<='Z';
					WHEN	1259	=>	bit_input<='Z';
					WHEN	1260	=>	bit_input<='Z';
					WHEN	1261	=>	bit_input<='Z';
					WHEN	1262	=>	bit_input<='Z';
					WHEN	1263	=>	bit_input<='Z';
					WHEN	1264	=>	bit_input<='Z';
					WHEN	1265	=>	bit_input<='Z';
					WHEN	1266	=>	bit_input<='Z';
					WHEN	1267	=>	bit_input<='Z';
					WHEN	1268	=>	bit_input<='Z';
					WHEN	1269	=>	bit_input<='Z';
					WHEN	1270	=>	bit_input<='Z';
					WHEN	1271	=>	bit_input<='Z';
					WHEN	1272	=>	bit_input<='Z';
					WHEN	1273	=>	bit_input<='Z';
					WHEN	1274	=>	bit_input<='Z';
					WHEN	1275	=>	bit_input<='Z';
					WHEN	1276	=>	bit_input<='Z';
					WHEN	1277	=>	bit_input<='Z';
					WHEN	1278	=>	bit_input<='Z';
					WHEN	1279	=>	bit_input<='Z';
					WHEN	1280	=>	bit_input<='Z';
					WHEN	1281	=>	bit_input<='Z';
					WHEN	1282	=>	bit_input<='Z';
					WHEN	1283	=>	bit_input<='Z';
					WHEN	1284	=>	bit_input<='Z';
					WHEN	1285	=>	bit_input<='Z';
					WHEN	1286	=>	bit_input<='Z';
					WHEN	1287	=>	bit_input<='Z';
					WHEN	1288	=>	bit_input<='Z';
					WHEN	1289	=>	bit_input<='Z';
					WHEN	1290	=>	bit_input<='Z';
					WHEN	1291	=>	bit_input<='Z';
					WHEN	1292	=>	bit_input<='Z';
					WHEN	1293	=>	bit_input<='Z';
					WHEN	1294	=>	bit_input<='Z';
					WHEN	1295	=>	bit_input<='Z';
					WHEN	1296	=>	bit_input<='Z';
					WHEN	1297	=>	bit_input<='Z';
					WHEN	1298	=>	bit_input<='Z';
					WHEN	1299	=>	bit_input<='Z';
					WHEN	1300	=>	bit_input<='Z';
					WHEN	1301	=>	bit_input<='Z';
					WHEN	1302	=>	bit_input<='Z';
					WHEN	1303	=>	bit_input<='Z';
					WHEN	1304	=>	bit_input<='Z';
					WHEN	1305	=>	bit_input<='Z';
					WHEN	1306	=>	bit_input<='Z';
					WHEN	1307	=>	bit_input<='Z';
					WHEN	1308	=>	bit_input<='Z';
					WHEN	1309	=>	bit_input<='Z';
					WHEN	1310	=>	bit_input<='Z';
					WHEN	1311	=>	bit_input<='Z';
					WHEN	1312	=>	bit_input<='Z';
					WHEN	1313	=>	bit_input<='Z';
					WHEN	1314	=>	bit_input<='Z';
					WHEN	1315	=>	bit_input<='Z';
					WHEN	1316	=>	bit_input<='Z';
					WHEN	1317	=>	bit_input<='Z';
					WHEN	1318	=>	bit_input<='Z';
					WHEN	1319	=>	bit_input<='Z';
					WHEN	1320	=>	bit_input<='Z';
					WHEN	1321	=>	bit_input<='Z';
					WHEN	1322	=>	bit_input<='Z';
					WHEN	1323	=>	bit_input<='Z';
					WHEN	1324	=>	bit_input<='Z';
					WHEN	1325	=>	bit_input<='Z';
					WHEN	1326	=>	bit_input<='Z';
					WHEN	1327	=>	bit_input<='Z';
					WHEN	1328	=>	bit_input<='Z';
					WHEN	1329	=>	bit_input<='Z';
					WHEN	1330	=>	bit_input<='Z';
					WHEN	1331	=>	bit_input<='Z';
					WHEN	1332	=>	bit_input<='Z';
					WHEN	1333	=>	bit_input<='Z';
					WHEN	1334	=>	bit_input<='Z';
					WHEN	1335	=>	bit_input<='Z';
					WHEN	1336	=>	bit_input<='Z';
					WHEN	1337	=>	bit_input<='Z';
					WHEN	1338	=>	bit_input<='Z';
					WHEN	1339	=>	bit_input<='Z';
					WHEN	1340	=>	bit_input<='Z';
					WHEN	1341	=>	bit_input<='Z';
					WHEN	1342	=>	bit_input<='Z';
					WHEN	1343	=>	bit_input<='Z';
					WHEN	1344	=>	bit_input<='Z';
					WHEN	1345	=>	bit_input<='Z';
					WHEN	1346	=>	bit_input<='Z';
					WHEN	1347	=>	bit_input<='Z';
					WHEN	1348	=>	bit_input<='Z';
					WHEN	1349	=>	bit_input<='Z';
					WHEN	1350	=>	bit_input<='Z';
					WHEN	1351	=>	bit_input<='Z';
					WHEN	1352	=>	bit_input<='Z';
					WHEN	1353	=>	bit_input<='Z';
					WHEN	1354	=>	bit_input<='Z';
					WHEN	1355	=>	bit_input<='Z';
					WHEN	1356	=>	bit_input<='Z';
					WHEN	1357	=>	bit_input<='Z';
					WHEN	1358	=>	bit_input<='Z';
					WHEN	1359	=>	bit_input<='Z';
					WHEN	1360	=>	bit_input<='Z';
					WHEN	1361	=>	bit_input<='Z';
					WHEN	1362	=>	bit_input<='Z';
					WHEN	1363	=>	bit_input<='Z';
					WHEN	1364	=>	bit_input<='Z';
					WHEN	1365	=>	bit_input<='Z';
					WHEN	1366	=>	bit_input<='Z';
					WHEN	1367	=>	bit_input<='Z';
					WHEN	1368	=>	bit_input<='Z';
					WHEN	1369	=>	bit_input<='Z';
					WHEN	1370	=>	bit_input<='Z';
					WHEN	1371	=>	bit_input<='Z';
					WHEN	1372	=>	bit_input<='Z';
					WHEN	1373	=>	bit_input<='Z';
					WHEN	1374	=>	bit_input<='Z';
					WHEN	1375	=>	bit_input<='Z';
					WHEN	1376	=>	bit_input<='Z';
					WHEN	1377	=>	bit_input<='Z';
					WHEN	1378	=>	bit_input<='Z';
					WHEN	1379	=>	bit_input<='Z';
					WHEN	1380	=>	bit_input<='Z';
					WHEN	1381	=>	bit_input<='Z';
					WHEN	1382	=>	bit_input<='Z';
					WHEN	1383	=>	bit_input<='Z';
					WHEN	1384	=>	bit_input<='Z';
					WHEN	1385	=>	bit_input<='Z';
					WHEN	1386	=>	bit_input<='Z';
					WHEN	1387	=>	bit_input<='Z';
					WHEN	1388	=>	bit_input<='Z';
					WHEN	1389	=>	bit_input<='Z';
					WHEN	1390	=>	bit_input<='Z';
					WHEN	1391	=>	bit_input<='Z';
					WHEN	1392	=>	bit_input<='Z';
					WHEN	1393	=>	bit_input<='Z';
					WHEN	1394	=>	bit_input<='Z';
					WHEN	1395	=>	bit_input<='Z';
					WHEN	1396	=>	bit_input<='Z';
					WHEN	1397	=>	bit_input<='Z';
					WHEN	1398	=>	bit_input<='Z';
					WHEN	1399	=>	bit_input<='Z';
					WHEN	1400	=>	bit_input<='Z';
					WHEN	1401	=>	bit_input<='Z';
					WHEN	1402	=>	bit_input<='Z';
					WHEN	1403	=>	bit_input<='Z';
					WHEN	1404	=>	bit_input<='Z';
					WHEN	1405	=>	bit_input<='Z';
					WHEN	1406	=>	bit_input<='Z';
					WHEN	1407	=>	bit_input<='Z';
					WHEN	1408	=>	bit_input<='Z';
					WHEN	1409	=>	bit_input<='Z';
					WHEN	1410	=>	bit_input<='Z';
					WHEN	1411	=>	bit_input<='Z';
					WHEN	1412	=>	bit_input<='Z';
					WHEN	1413	=>	bit_input<='Z';
					WHEN	1414	=>	bit_input<='Z';
					WHEN	1415	=>	bit_input<='Z';
					WHEN	1416	=>	bit_input<='Z';
					WHEN	1417	=>	bit_input<='Z';
					WHEN	1418	=>	bit_input<='Z';
					WHEN	1419	=>	bit_input<='Z';
					WHEN	1420	=>	bit_input<='Z';
					WHEN	1421	=>	bit_input<='Z';
					WHEN	1422	=>	bit_input<='Z';
					WHEN	1423	=>	bit_input<='Z';
					WHEN	1424	=>	bit_input<='Z';
					WHEN	1425	=>	bit_input<='Z';
					WHEN	1426	=>	bit_input<='Z';
					WHEN	1427	=>	bit_input<='Z';
					WHEN	1428	=>	bit_input<='Z';
					WHEN	1429	=>	bit_input<='Z';
					WHEN	1430	=>	bit_input<='Z';
					WHEN	1431	=>	bit_input<='Z';
					WHEN	1432	=>	bit_input<='Z';
					WHEN	1433	=>	bit_input<='Z';
					WHEN	1434	=>	bit_input<='Z';
					WHEN	1435	=>	bit_input<='Z';
					WHEN	1436	=>	bit_input<='Z';
					WHEN	1437	=>	bit_input<='Z';
					WHEN	1438	=>	bit_input<='Z';
					WHEN	1439	=>	bit_input<='Z';
					WHEN	1440	=>	bit_input<='Z';
					WHEN	1441	=>	bit_input<='Z';
					WHEN	1442	=>	bit_input<='Z';
					WHEN	1443	=>	bit_input<='Z';
					WHEN	1444	=>	bit_input<='Z';
					WHEN	1445	=>	bit_input<='Z';
					WHEN	1446	=>	bit_input<='Z';
					WHEN	1447	=>	bit_input<='Z';
					WHEN	1448	=>	bit_input<='Z';
					WHEN	1449	=>	bit_input<='Z';
					WHEN	1450	=>	bit_input<='Z';
					WHEN	1451	=>	bit_input<='Z';
					WHEN	1452	=>	bit_input<='Z';
					WHEN	1453	=>	bit_input<='Z';
					WHEN	1454	=>	bit_input<='Z';
					WHEN	1455	=>	bit_input<='Z';
					WHEN	1456	=>	bit_input<='Z';
					WHEN	1457	=>	bit_input<='Z';
					WHEN	1458	=>	bit_input<='Z';
					WHEN	1459	=>	bit_input<='Z';
					WHEN	1460	=>	bit_input<='Z';
					WHEN	1461	=>	bit_input<='Z';
					WHEN	1462	=>	bit_input<='Z';
					WHEN	1463	=>	bit_input<='Z';
					WHEN	1464	=>	bit_input<='Z';
					WHEN	1465	=>	bit_input<='Z';
					WHEN	1466	=>	bit_input<='Z';
					WHEN	1467	=>	bit_input<='Z';
					WHEN	1468	=>	bit_input<='Z';
					WHEN	1469	=>	bit_input<='Z';
					WHEN	1470	=>	bit_input<='Z';
					WHEN	1471	=>	bit_input<='Z';
					WHEN	1472	=>	bit_input<='Z';
					WHEN	1473	=>	bit_input<='Z';
					WHEN	1474	=>	bit_input<='Z';
					WHEN	1475	=>	bit_input<='Z';
					WHEN	1476	=>	bit_input<='Z';
					WHEN	1477	=>	bit_input<='Z';
					WHEN	1478	=>	bit_input<='Z';
					WHEN	1479	=>	bit_input<='Z';
					WHEN	1480	=>	bit_input<='Z';
					WHEN	1481	=>	bit_input<='Z';
					WHEN	1482	=>	bit_input<='Z';
					WHEN	1483	=>	bit_input<='Z';
					WHEN	1484	=>	bit_input<='Z';
					WHEN	1485	=>	bit_input<='Z';
					WHEN	1486	=>	bit_input<='Z';
					WHEN	1487	=>	bit_input<='Z';
					WHEN	1488	=>	bit_input<='Z';
					WHEN	1489	=>	bit_input<='Z';
					WHEN	1490	=>	bit_input<='Z';
					WHEN	1491	=>	bit_input<='Z';
					WHEN	1492	=>	bit_input<='Z';
					WHEN	1493	=>	bit_input<='Z';
					WHEN	1494	=>	bit_input<='Z';
					WHEN	1495	=>	bit_input<='Z';
					WHEN	1496	=>	bit_input<='Z';
					WHEN	1497	=>	bit_input<='Z';
					WHEN	1498	=>	bit_input<='Z';
					WHEN	1499	=>	bit_input<='Z';
					WHEN	1500	=>	bit_input<='Z';
					WHEN	1501	=>	bit_input<='Z';
					WHEN	1502	=>	bit_input<='Z';
					WHEN	1503	=>	bit_input<='Z';
					WHEN	1504	=>	bit_input<='Z';
					WHEN	1505	=>	bit_input<='Z';
					WHEN	1506	=>	bit_input<='Z';
					WHEN	1507	=>	bit_input<='Z';
					WHEN	1508	=>	bit_input<='Z';
					WHEN	1509	=>	bit_input<='Z';
					WHEN	1510	=>	bit_input<='Z';
					WHEN	1511	=>	bit_input<='Z';
					WHEN	1512	=>	bit_input<='Z';
					WHEN	1513	=>	bit_input<='Z';
					WHEN	1514	=>	bit_input<='Z';
					WHEN	1515	=>	bit_input<='Z';
					WHEN	1516	=>	bit_input<='Z';
					WHEN	1517	=>	bit_input<='Z';
					WHEN	1518	=>	bit_input<='Z';
					WHEN	1519	=>	bit_input<='Z';
					WHEN	1520	=>	bit_input<='Z';
					WHEN	1521	=>	bit_input<='Z';
					WHEN	1522	=>	bit_input<='Z';
					WHEN	1523	=>	bit_input<='Z';
					WHEN	1524	=>	bit_input<='Z';
					WHEN	1525	=>	bit_input<='Z';
					WHEN	1526	=>	bit_input<='Z';
					WHEN	1527	=>	bit_input<='Z';
					WHEN	1528	=>	bit_input<='Z';
					WHEN	1529	=>	bit_input<='Z';
					WHEN	1530	=>	bit_input<='Z';
					WHEN	1531	=>	bit_input<='Z';
					WHEN	1532	=>	bit_input<='Z';
					WHEN	1533	=>	bit_input<='Z';
					WHEN	1534	=>	bit_input<='Z';
					WHEN	1535	=>	bit_input<='Z';
					WHEN	1536	=>	bit_input<='Z';
					WHEN	1537	=>	bit_input<='Z';
					WHEN	1538	=>	bit_input<='Z';
					WHEN	1539	=>	bit_input<='Z';
					WHEN	1540	=>	bit_input<='Z';
					WHEN	1541	=>	bit_input<='Z';
					WHEN	1542	=>	bit_input<='Z';
					WHEN	1543	=>	bit_input<='Z';
					WHEN	1544	=>	bit_input<='Z';
					WHEN	1545	=>	bit_input<='Z';
					WHEN	1546	=>	bit_input<='Z';
					WHEN	1547	=>	bit_input<='Z';
					WHEN	1548	=>	bit_input<='Z';
					WHEN	1549	=>	bit_input<='Z';
					WHEN	1550	=>	bit_input<='Z';
					WHEN	1551	=>	bit_input<='Z';
					WHEN	1552	=>	bit_input<='Z';
					WHEN	1553	=>	bit_input<='Z';
					WHEN	1554	=>	bit_input<='Z';
					WHEN	1555	=>	bit_input<='Z';
					WHEN	1556	=>	bit_input<='Z';
					WHEN	1557	=>	bit_input<='Z';
					WHEN	1558	=>	bit_input<='Z';
					WHEN	1559	=>	bit_input<='Z';
					WHEN	1560	=>	bit_input<='Z';
					WHEN	1561	=>	bit_input<='Z';
					WHEN	1562	=>	bit_input<='Z';
					WHEN	1563	=>	bit_input<='Z';
					WHEN	1564	=>	bit_input<='Z';
					WHEN	1565	=>	bit_input<='Z';
					WHEN	1566	=>	bit_input<='Z';
					WHEN	1567	=>	bit_input<='Z';
					WHEN	1568	=>	bit_input<='Z';
					WHEN	1569	=>	bit_input<='Z';
					WHEN	1570	=>	bit_input<='Z';
					WHEN	1571	=>	bit_input<='Z';
					WHEN	1572	=>	bit_input<='Z';
					WHEN	1573	=>	bit_input<='Z';
					WHEN	1574	=>	bit_input<='Z';
					WHEN	1575	=>	bit_input<='Z';
					WHEN	1576	=>	bit_input<='Z';
					WHEN	1577	=>	bit_input<='Z';
					WHEN	1578	=>	bit_input<='Z';
					WHEN	1579	=>	bit_input<='Z';
					WHEN	1580	=>	bit_input<='Z';
					WHEN	1581	=>	bit_input<='Z';
					WHEN	1582	=>	bit_input<='Z';
					WHEN	1583	=>	bit_input<='Z';
					WHEN	1584	=>	bit_input<='Z';
					WHEN	1585	=>	bit_input<='Z';
					WHEN	1586	=>	bit_input<='Z';
					WHEN	1587	=>	bit_input<='Z';
					WHEN	1588	=>	bit_input<='Z';
					WHEN	1589	=>	bit_input<='Z';
					WHEN	1590	=>	bit_input<='Z';
					WHEN	1591	=>	bit_input<='Z';
					WHEN	1592	=>	bit_input<='Z';
					WHEN	1593	=>	bit_input<='Z';
					WHEN	1594	=>	bit_input<='Z';
					WHEN	1595	=>	bit_input<='Z';
					WHEN	1596	=>	bit_input<='Z';
					WHEN	1597	=>	bit_input<='Z';
					WHEN	1598	=>	bit_input<='Z';
					WHEN	1599	=>	bit_input<='Z';
					WHEN	1600	=>	bit_input<='Z';
					WHEN	1601	=>	bit_input<='Z';
					WHEN	1602	=>	bit_input<='Z';
					WHEN	1603	=>	bit_input<='Z';
					WHEN	1604	=>	bit_input<='Z';
					WHEN	1605	=>	bit_input<='Z';
					WHEN	1606	=>	bit_input<='Z';
					WHEN	1607	=>	bit_input<='Z';
					WHEN	1608	=>	bit_input<='Z';
					WHEN	1609	=>	bit_input<='Z';
					WHEN	1610	=>	bit_input<='Z';
					WHEN	1611	=>	bit_input<='Z';
					WHEN	1612	=>	bit_input<='Z';
					WHEN	1613	=>	bit_input<='Z';
					WHEN	1614	=>	bit_input<='Z';
					WHEN	1615	=>	bit_input<='Z';
					WHEN	1616	=>	bit_input<='Z';
					WHEN	1617	=>	bit_input<='Z';
					WHEN	1618	=>	bit_input<='Z';
					WHEN	1619	=>	bit_input<='Z';
					WHEN	1620	=>	bit_input<='Z';
					WHEN	1621	=>	bit_input<='Z';
					WHEN	1622	=>	bit_input<='Z';
					WHEN	1623	=>	bit_input<='Z';
					WHEN	1624	=>	bit_input<='Z';
					WHEN	1625	=>	bit_input<='Z';
					WHEN	1626	=>	bit_input<='Z';
					WHEN	1627	=>	bit_input<='Z';
					WHEN	1628	=>	bit_input<='Z';
					WHEN	1629	=>	bit_input<='Z';
					WHEN	1630	=>	bit_input<='Z';
					WHEN	1631	=>	bit_input<='Z';
					WHEN	1632	=>	bit_input<='Z';
					WHEN	1633	=>	bit_input<='Z';
					WHEN	1634	=>	bit_input<='Z';
					WHEN	1635	=>	bit_input<='Z';
					WHEN	1636	=>	bit_input<='Z';
					WHEN	1637	=>	bit_input<='Z';
					WHEN	1638	=>	bit_input<='Z';
					WHEN	1639	=>	bit_input<='Z';
					WHEN	1640	=>	bit_input<='Z';
					WHEN	1641	=>	bit_input<='Z';
					WHEN	1642	=>	bit_input<='Z';
					WHEN	1643	=>	bit_input<='Z';
					WHEN	1644	=>	bit_input<='Z';
					WHEN	1645	=>	bit_input<='Z';
					WHEN	1646	=>	bit_input<='Z';
					WHEN	1647	=>	bit_input<='Z';
					WHEN	1648	=>	bit_input<='Z';
					WHEN	1649	=>	bit_input<='Z';
					WHEN	1650	=>	bit_input<='Z';
					WHEN	1651	=>	bit_input<='Z';
					WHEN	1652	=>	bit_input<='Z';
					WHEN	1653	=>	bit_input<='Z';
					WHEN	1654	=>	bit_input<='Z';
					WHEN	1655	=>	bit_input<='Z';
					WHEN	1656	=>	bit_input<='Z';
					WHEN	1657	=>	bit_input<='Z';
					WHEN	1658	=>	bit_input<='Z';
					WHEN	1659	=>	bit_input<='Z';
					WHEN	1660	=>	bit_input<='Z';
					WHEN	1661	=>	bit_input<='Z';
					WHEN	1662	=>	bit_input<='Z';
					WHEN	1663	=>	bit_input<='Z';
					WHEN	1664	=>	bit_input<='Z';
					WHEN	1665	=>	bit_input<='Z';
					WHEN	1666	=>	bit_input<='Z';
					WHEN	1667	=>	bit_input<='Z';
					WHEN	1668	=>	bit_input<='Z';
					WHEN	1669	=>	bit_input<='Z';
					WHEN	1670	=>	bit_input<='Z';
					WHEN	1671	=>	bit_input<='Z';
					WHEN	1672	=>	bit_input<='Z';
					WHEN	1673	=>	bit_input<='Z';
					WHEN	1674	=>	bit_input<='Z';
					WHEN	1675	=>	bit_input<='Z';
					WHEN	1676	=>	bit_input<='Z';
					WHEN	1677	=>	bit_input<='Z';
					WHEN	1678	=>	bit_input<='Z';
					WHEN	1679	=>	bit_input<='Z';
					WHEN	1680	=>	bit_input<='Z';
					WHEN	1681	=>	bit_input<='Z';
					WHEN	1682	=>	bit_input<='Z';
					WHEN	1683	=>	bit_input<='Z';
					WHEN	1684	=>	bit_input<='Z';
					WHEN	1685	=>	bit_input<='Z';
					WHEN	1686	=>	bit_input<='Z';
					WHEN	1687	=>	bit_input<='Z';
					WHEN	1688	=>	bit_input<='Z';
					WHEN	1689	=>	bit_input<='Z';
					WHEN	1690	=>	bit_input<='Z';
					WHEN	1691	=>	bit_input<='Z';
					WHEN	1692	=>	bit_input<='Z';
					WHEN	1693	=>	bit_input<='Z';
					WHEN	1694	=>	bit_input<='Z';
					WHEN	1695	=>	bit_input<='Z';
					WHEN	1696	=>	bit_input<='Z';
					WHEN	1697	=>	bit_input<='Z';
					WHEN	1698	=>	bit_input<='Z';
					WHEN	1699	=>	bit_input<='Z';
					WHEN	1700	=>	bit_input<='Z';
					WHEN	1701	=>	bit_input<='Z';
					WHEN	1702	=>	bit_input<='Z';
					WHEN	1703	=>	bit_input<='Z';
					WHEN	1704	=>	bit_input<='Z';
					WHEN	1705	=>	bit_input<='Z';
					WHEN	1706	=>	bit_input<='Z';
					WHEN	1707	=>	bit_input<='Z';
					WHEN	1708	=>	bit_input<='Z';
					WHEN	1709	=>	bit_input<='Z';
					WHEN	1710	=>	bit_input<='Z';
					WHEN	1711	=>	bit_input<='Z';
					WHEN	1712	=>	bit_input<='Z';
					WHEN	1713	=>	bit_input<='Z';
					WHEN	1714	=>	bit_input<='Z';
					WHEN	1715	=>	bit_input<='Z';
					WHEN	1716	=>	bit_input<='Z';
					WHEN	1717	=>	bit_input<='Z';
					WHEN	1718	=>	bit_input<='Z';
					WHEN	1719	=>	bit_input<='Z';
					WHEN	1720	=>	bit_input<='Z';
					WHEN	1721	=>	bit_input<='Z';
					WHEN	1722	=>	bit_input<='Z';
					WHEN	1723	=>	bit_input<='Z';
					WHEN	1724	=>	bit_input<='Z';
					WHEN	1725	=>	bit_input<='Z';
					WHEN	1726	=>	bit_input<='Z';
					WHEN	1727	=>	bit_input<='Z';
					WHEN	1728	=>	bit_input<='Z';
					WHEN	1729	=>	bit_input<='Z';
					WHEN	1730	=>	bit_input<='Z';
					WHEN	1731	=>	bit_input<='Z';
					WHEN	1732	=>	bit_input<='Z';
					WHEN	1733	=>	bit_input<='Z';
					WHEN	1734	=>	bit_input<='Z';
					WHEN	1735	=>	bit_input<='Z';
					WHEN	1736	=>	bit_input<='Z';
					WHEN	1737	=>	bit_input<='Z';
					WHEN	1738	=>	bit_input<='Z';
					WHEN	1739	=>	bit_input<='Z';
					WHEN	1740	=>	bit_input<='Z';
					WHEN	1741	=>	bit_input<='Z';
					WHEN	1742	=>	bit_input<='Z';
					WHEN	1743	=>	bit_input<='Z';
					WHEN	1744	=>	bit_input<='Z';
					WHEN	1745	=>	bit_input<='Z';
					WHEN	1746	=>	bit_input<='Z';
					WHEN	1747	=>	bit_input<='Z';
					WHEN	1748	=>	bit_input<='Z';
					WHEN	1749	=>	bit_input<='Z';
					WHEN	1750	=>	bit_input<='Z';
					WHEN	1751	=>	bit_input<='Z';
					WHEN	1752	=>	bit_input<='Z';
					WHEN	1753	=>	bit_input<='Z';
					WHEN	1754	=>	bit_input<='Z';
					WHEN	1755	=>	bit_input<='Z';
					WHEN	1756	=>	bit_input<='Z';
					WHEN	1757	=>	bit_input<='Z';
					WHEN	1758	=>	bit_input<='Z';
					WHEN	1759	=>	bit_input<='Z';
					WHEN	1760	=>	bit_input<='Z';
					WHEN	1761	=>	bit_input<='Z';
					WHEN	1762	=>	bit_input<='Z';
					WHEN	1763	=>	bit_input<='Z';
					WHEN	1764	=>	bit_input<='Z';
					WHEN	1765	=>	bit_input<='Z';
					WHEN	1766	=>	bit_input<='Z';
					WHEN	1767	=>	bit_input<='Z';
					WHEN	1768	=>	bit_input<='Z';
					WHEN	1769	=>	bit_input<='Z';
					WHEN	1770	=>	bit_input<='Z';
					WHEN	1771	=>	bit_input<='Z';
					WHEN	1772	=>	bit_input<='Z';
					WHEN	1773	=>	bit_input<='Z';
					WHEN	1774	=>	bit_input<='Z';
					WHEN	1775	=>	bit_input<='Z';
					WHEN	1776	=>	bit_input<='Z';
					WHEN	1777	=>	bit_input<='Z';
					WHEN	1778	=>	bit_input<='Z';
					WHEN	1779	=>	bit_input<='Z';
					WHEN	1780	=>	bit_input<='Z';
					WHEN	1781	=>	bit_input<='Z';
					WHEN	1782	=>	bit_input<='Z';
					WHEN	1783	=>	bit_input<='Z';
					WHEN	1784	=>	bit_input<='Z';
					WHEN	1785	=>	bit_input<='Z';
					WHEN	1786	=>	bit_input<='Z';
					WHEN	1787	=>	bit_input<='Z';
					WHEN	1788	=>	bit_input<='Z';
					WHEN	1789	=>	bit_input<='Z';
					WHEN	1790	=>	bit_input<='Z';
					WHEN	1791	=>	bit_input<='Z';
					WHEN	1792	=>	bit_input<='Z';
					WHEN	1793	=>	bit_input<='Z';
					WHEN	1794	=>	bit_input<='Z';
					WHEN	1795	=>	bit_input<='Z';
					WHEN	1796	=>	bit_input<='Z';
					WHEN	1797	=>	bit_input<='Z';
					WHEN	1798	=>	bit_input<='Z';
					WHEN	1799	=>	bit_input<='Z';
					WHEN	1800	=>	bit_input<='Z';
					WHEN	1801	=>	bit_input<='Z';
					WHEN	1802	=>	bit_input<='Z';
					WHEN	1803	=>	bit_input<='Z';
					WHEN	1804	=>	bit_input<='Z';
					WHEN	1805	=>	bit_input<='Z';
					WHEN	1806	=>	bit_input<='Z';
					WHEN	1807	=>	bit_input<='Z';
					WHEN	1808	=>	bit_input<='Z';
					WHEN	1809	=>	bit_input<='Z';
					WHEN	1810	=>	bit_input<='Z';
					WHEN	1811	=>	bit_input<='Z';
					WHEN	1812	=>	bit_input<='Z';
					WHEN	1813	=>	bit_input<='Z';
					WHEN	1814	=>	bit_input<='Z';
					WHEN	1815	=>	bit_input<='Z';
					WHEN	1816	=>	bit_input<='Z';
					WHEN	1817	=>	bit_input<='Z';
					WHEN	1818	=>	bit_input<='Z';
					WHEN	1819	=>	bit_input<='Z';
					WHEN	1820	=>	bit_input<='Z';
					WHEN	1821	=>	bit_input<='Z';
					WHEN	1822	=>	bit_input<='Z';
					WHEN	1823	=>	bit_input<='Z';
					WHEN	1824	=>	bit_input<='Z';
					WHEN	1825	=>	bit_input<='Z';
					WHEN	1826	=>	bit_input<='Z';
					WHEN	1827	=>	bit_input<='Z';
					WHEN	1828	=>	bit_input<='Z';
					WHEN	1829	=>	bit_input<='Z';
					WHEN	1830	=>	bit_input<='Z';
					WHEN	1831	=>	bit_input<='Z';
					WHEN	1832	=>	bit_input<='Z';
					WHEN	1833	=>	bit_input<='Z';
					WHEN	1834	=>	bit_input<='Z';
					WHEN	1835	=>	bit_input<='Z';
					WHEN	1836	=>	bit_input<='Z';
					WHEN	1837	=>	bit_input<='Z';
					WHEN	1838	=>	bit_input<='Z';
					WHEN	1839	=>	bit_input<='Z';
					WHEN	1840	=>	bit_input<='Z';
					WHEN	1841	=>	bit_input<='Z';
					WHEN	1842	=>	bit_input<='Z';
					WHEN	1843	=>	bit_input<='Z';
					WHEN	1844	=>	bit_input<='Z';
					WHEN	1845	=>	bit_input<='Z';
					WHEN	1846	=>	bit_input<='Z';
					WHEN	1847	=>	bit_input<='Z';
					WHEN	1848	=>	bit_input<='Z';
					WHEN	1849	=>	bit_input<='Z';
					WHEN	1850	=>	bit_input<='Z';
					WHEN	1851	=>	bit_input<='Z';
					WHEN	1852	=>	bit_input<='Z';
					WHEN	1853	=>	bit_input<='Z';
					WHEN	1854	=>	bit_input<='Z';
					WHEN	1855	=>	bit_input<='Z';
					WHEN	1856	=>	bit_input<='Z';
					WHEN	1857	=>	bit_input<='Z';
					WHEN	1858	=>	bit_input<='Z';
					WHEN	1859	=>	bit_input<='Z';
					WHEN	1860	=>	bit_input<='Z';
					WHEN	1861	=>	bit_input<='Z';
					WHEN	1862	=>	bit_input<='Z';
					WHEN	1863	=>	bit_input<='Z';
					WHEN	1864	=>	bit_input<='Z';
					WHEN	1865	=>	bit_input<='Z';
					WHEN	1866	=>	bit_input<='Z';
					WHEN	1867	=>	bit_input<='Z';
					WHEN	1868	=>	bit_input<='Z';
					WHEN	1869	=>	bit_input<='Z';
					WHEN	1870	=>	bit_input<='Z';
					WHEN	1871	=>	bit_input<='Z';
					WHEN	1872	=>	bit_input<='Z';
					WHEN	1873	=>	bit_input<='Z';
					WHEN	1874	=>	bit_input<='Z';
					WHEN	1875	=>	bit_input<='Z';
					WHEN	1876	=>	bit_input<='Z';
					WHEN	1877	=>	bit_input<='Z';
					WHEN	1878	=>	bit_input<='Z';
					WHEN	1879	=>	bit_input<='Z';
					WHEN	1880	=>	bit_input<='Z';
					WHEN	1881	=>	bit_input<='Z';
					WHEN	1882	=>	bit_input<='Z';
					WHEN	1883	=>	bit_input<='Z';
					WHEN	1884	=>	bit_input<='Z';
					WHEN	1885	=>	bit_input<='Z';
					WHEN	1886	=>	bit_input<='Z';
					WHEN	1887	=>	bit_input<='Z';
					WHEN	1888	=>	bit_input<='Z';
					WHEN	1889	=>	bit_input<='Z';
					WHEN	1890	=>	bit_input<='Z';
					WHEN	1891	=>	bit_input<='Z';
					WHEN	1892	=>	bit_input<='Z';
					WHEN	1893	=>	bit_input<='Z';
					WHEN	1894	=>	bit_input<='Z';
					WHEN	1895	=>	bit_input<='Z';
					WHEN	1896	=>	bit_input<='Z';
					WHEN	1897	=>	bit_input<='Z';
					WHEN	1898	=>	bit_input<='Z';
					WHEN	1899	=>	bit_input<='Z';
					WHEN	1900	=>	bit_input<='Z';
					WHEN	1901	=>	bit_input<='Z';
					WHEN	1902	=>	bit_input<='Z';
					WHEN	1903	=>	bit_input<='Z';
					WHEN	1904	=>	bit_input<='Z';
					WHEN	1905	=>	bit_input<='Z';
					WHEN	1906	=>	bit_input<='Z';
					WHEN	1907	=>	bit_input<='Z';
					WHEN	1908	=>	bit_input<='Z';
					WHEN	1909	=>	bit_input<='Z';
					WHEN	1910	=>	bit_input<='Z';
					WHEN	1911	=>	bit_input<='Z';
					WHEN	1912	=>	bit_input<='Z';
					WHEN	1913	=>	bit_input<='Z';
					WHEN	1914	=>	bit_input<='Z';
					WHEN	1915	=>	bit_input<='Z';
					WHEN	1916	=>	bit_input<='Z';
					WHEN	1917	=>	bit_input<='Z';
					WHEN	1918	=>	bit_input<='Z';
					WHEN	1919	=>	bit_input<='Z';
					WHEN	1920	=>	bit_input<='Z';
					WHEN	1921	=>	bit_input<='Z';
					WHEN	1922	=>	bit_input<='Z';
					WHEN	1923	=>	bit_input<='Z';
					WHEN	1924	=>	bit_input<='Z';
					WHEN	1925	=>	bit_input<='Z';
					WHEN	1926	=>	bit_input<='Z';
					WHEN	1927	=>	bit_input<='Z';
					WHEN	1928	=>	bit_input<='Z';
					WHEN	1929	=>	bit_input<='Z';
					WHEN	1930	=>	bit_input<='Z';
					WHEN	1931	=>	bit_input<='Z';
					WHEN	1932	=>	bit_input<='Z';
					WHEN	1933	=>	bit_input<='Z';
					WHEN	1934	=>	bit_input<='Z';
					WHEN	1935	=>	bit_input<='Z';
					WHEN	1936	=>	bit_input<='Z';
					WHEN	1937	=>	bit_input<='Z';
					WHEN	1938	=>	bit_input<='Z';
					WHEN	1939	=>	bit_input<='Z';
					WHEN	1940	=>	bit_input<='Z';
					WHEN	1941	=>	bit_input<='Z';
					WHEN	1942	=>	bit_input<='Z';
					WHEN	1943	=>	bit_input<='Z';
					WHEN	1944	=>	bit_input<='Z';
					WHEN	1945	=>	bit_input<='Z';
					WHEN	1946	=>	bit_input<='Z';
					WHEN	1947	=>	bit_input<='Z';
					WHEN	1948	=>	bit_input<='Z';
					WHEN	1949	=>	bit_input<='Z';
					WHEN	1950	=>	bit_input<='Z';
					WHEN	1951	=>	bit_input<='Z';
					WHEN	1952	=>	bit_input<='Z';
					WHEN	1953	=>	bit_input<='Z';
					WHEN	1954	=>	bit_input<='Z';
					WHEN	1955	=>	bit_input<='Z';
					WHEN	1956	=>	bit_input<='Z';
					WHEN	1957	=>	bit_input<='Z';
					WHEN	1958	=>	bit_input<='Z';
					WHEN	1959	=>	bit_input<='Z';
					WHEN	1960	=>	bit_input<='Z';
					WHEN	1961	=>	bit_input<='Z';
					WHEN	1962	=>	bit_input<='Z';
					WHEN	1963	=>	bit_input<='Z';
					WHEN	1964	=>	bit_input<='Z';
					WHEN	1965	=>	bit_input<='Z';
					WHEN	1966	=>	bit_input<='Z';
					WHEN	1967	=>	bit_input<='Z';
					WHEN	1968	=>	bit_input<='Z';
					WHEN	1969	=>	bit_input<='Z';
					WHEN	1970	=>	bit_input<='Z';
					WHEN	1971	=>	bit_input<='Z';
					WHEN	1972	=>	bit_input<='Z';
					WHEN	1973	=>	bit_input<='Z';
					WHEN	1974	=>	bit_input<='Z';
					WHEN	1975	=>	bit_input<='Z';
					WHEN	1976	=>	bit_input<='Z';
					WHEN	1977	=>	bit_input<='Z';
					WHEN	1978	=>	bit_input<='Z';
					WHEN	1979	=>	bit_input<='Z';
					WHEN	1980	=>	bit_input<='Z';
					WHEN	1981	=>	bit_input<='Z';
					WHEN	1982	=>	bit_input<='Z';
					WHEN	1983	=>	bit_input<='Z';
					WHEN	1984	=>	bit_input<='Z';
					WHEN	1985	=>	bit_input<='Z';
					WHEN	1986	=>	bit_input<='Z';
					WHEN	1987	=>	bit_input<='Z';
					WHEN	1988	=>	bit_input<='Z';
					WHEN	1989	=>	bit_input<='Z';
					WHEN	1990	=>	bit_input<='Z';
					WHEN	1991	=>	bit_input<='Z';
					WHEN	1992	=>	bit_input<='Z';
					WHEN	1993	=>	bit_input<='Z';
					WHEN	1994	=>	bit_input<='Z';
					WHEN	1995	=>	bit_input<='Z';
					WHEN	1996	=>	bit_input<='Z';
					WHEN	1997	=>	bit_input<='Z';
					WHEN	1998	=>	bit_input<='Z';
					WHEN	1999	=>	bit_input<='Z';
					WHEN	2000	=>	bit_input<='Z';
					WHEN	2001	=>	bit_input<='Z';
					WHEN	2002	=>	bit_input<='Z';
					WHEN	2003	=>	bit_input<='Z';
					WHEN	2004	=>	bit_input<='Z';
					WHEN	2005	=>	bit_input<='Z';
					WHEN	2006	=>	bit_input<='Z';
					WHEN	2007	=>	bit_input<='Z';
					WHEN	2008	=>	bit_input<='Z';
					WHEN	2009	=>	bit_input<='Z';
					WHEN	2010	=>	bit_input<='Z';
					WHEN	2011	=>	bit_input<='Z';
					WHEN	2012	=>	bit_input<='Z';
					WHEN	2013	=>	bit_input<='Z';
					WHEN	2014	=>	bit_input<='Z';
					WHEN	2015	=>	bit_input<='Z';
					WHEN	2016	=>	bit_input<='Z';
					WHEN	2017	=>	bit_input<='Z';
					WHEN	2018	=>	bit_input<='Z';
					WHEN	2019	=>	bit_input<='Z';
					WHEN	2020	=>	bit_input<='Z';
					WHEN	2021	=>	bit_input<='Z';
					WHEN	2022	=>	bit_input<='Z';
					WHEN	2023	=>	bit_input<='Z';
					WHEN	2024	=>	bit_input<='Z';
					WHEN	2025	=>	bit_input<='Z';
					WHEN	2026	=>	bit_input<='Z';
					WHEN	2027	=>	bit_input<='Z';
					WHEN	2028	=>	bit_input<='Z';
					WHEN	2029	=>	bit_input<='Z';
					WHEN	2030	=>	bit_input<='Z';
					WHEN	2031	=>	bit_input<='Z';
					WHEN	2032	=>	bit_input<='Z';
					WHEN	2033	=>	bit_input<='Z';
					WHEN	2034	=>	bit_input<='Z';
					WHEN	2035	=>	bit_input<='Z';
					WHEN	2036	=>	bit_input<='Z';
					WHEN	2037	=>	bit_input<='Z';
					WHEN	2038	=>	bit_input<='Z';
					WHEN	2039	=>	bit_input<='Z';
					WHEN	2040	=>	bit_input<='Z';
					WHEN	2041	=>	bit_input<='Z';
					WHEN	2042	=>	bit_input<='Z';
					WHEN	2043	=>	bit_input<='Z';
					WHEN	2044	=>	bit_input<='Z';
					WHEN	2045	=>	bit_input<='Z';
					WHEN	2046	=>	bit_input<='Z';
					WHEN	2047	=>	bit_input<='Z';
					WHEN	2048	=>	bit_input<='Z';
					WHEN	len 	=>	testing<=False;
					WHEN	OTHERS	=>	NULL;
				END CASE;
				if clock = '1' and clock'event then 
					count:= count + 1;
				END IF;

		END PROCESS proc_test;
END interleaver_test_arch;